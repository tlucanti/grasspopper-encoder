`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////
// Company: Miet
// Engineer: Kostya
// 
// Create Date: 19.06.2022 13:07:40
// Design Name: Grasspopper
// Module Name: non_linear
// Project Name: Grasspopper
// Target Devices: any
// Tool Versions: 2021.1
// Description:
//   sync module
//   module implements non_linear action in one stage for grasspopper encoding
//
// Parameters:
//   rst            - reset signal
//   clk            - clock signal
//   data_i         - 255 bit (16 bytes) data to be encoded
//   data_o         - 255 bit (16 bytes) encoded data
//
// Dependencies: None
// 
// Revision: v0.1
//   v0.1 - file Created
//
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module non_linear(data_i, data_o);

input [127:0]   data_i;
/*

*/

output [127:0]  data_o;
/*

*/

wire [7:0] extra_byte;
wire [7:0] extra_byte_0;
wire [7:0] extra_byte_1;
wire [7:0] extra_byte_2;
wire [7:0] extra_byte_3;
wire [7:0] extra_byte_4;
wire [7:0] extra_byte_5;
wire [7:0] extra_byte_6;
wire [7:0] extra_byte_7;
wire [7:0] extra_byte_8;
wire [7:0] extra_byte_9;
wire [7:0] extra_byte_A;
wire [7:0] extra_byte_B;
wire [7:0] extra_byte_C;
wire [7:0] extra_byte_D;
wire [7:0] extra_byte_E;
wire [7:0] extra_byte_F;

assign extra_byte = 
    extra_byte_0 ^
    extra_byte_1 ^
    extra_byte_2 ^
    extra_byte_3 ^
    extra_byte_4 ^
    extra_byte_5 ^
    extra_byte_6 ^
    extra_byte_7 ^
    extra_byte_8 ^
    extra_byte_9 ^
    extra_byte_A ^
    extra_byte_B ^
    extra_byte_C ^
    extra_byte_D ^
    extra_byte_E ^
    extra_byte_F;

assign extra_byte_0 =    galois_lookup_148(data_i[127:120]);
assign extra_byte_1 =    galois_lookup_032(data_i[119:112]);
assign extra_byte_2 =    galois_lookup_133(data_i[111:104]);
assign extra_byte_3 =    galois_lookup_016(data_i[103:096]);
assign extra_byte_4 =    galois_lookup_194(data_i[095:088]);
assign extra_byte_5 =    galois_lookup_192(data_i[087:080]);
assign extra_byte_6 =                      data_i[079:072] ;
assign extra_byte_7 =    galois_lookup_251(data_i[071:064]);
assign extra_byte_8 =                      data_i[063:056] ;
assign extra_byte_9 =    galois_lookup_192(data_i[055:048]);
assign extra_byte_B =    galois_lookup_194(data_i[047:040]);
assign extra_byte_A =    galois_lookup_016(data_i[039:032]);
assign extra_byte_C =    galois_lookup_133(data_i[031:024]);
assign extra_byte_D =    galois_lookup_032(data_i[023:016]);
assign extra_byte_E =    galois_lookup_148(data_i[015:008]);
assign extra_byte_F =                      data_i[007:000] ;

assign data_o = {extra_byte, data_i[127:008]};

// -----------------------------------------------------------------------------
function automatic [7:0] xor_reduce;
/*

*/
    input   [127:0] data;

    begin
        xor_reduce =    data[015:008] ^ data[023:016] ^ data[031:024] ^
                        data[039:032] ^ data[047:040] ^ data[055:048] ^
                        data[063:056] ^ data[071:064] ^ data[079:072] ^
                        data[087:080] ^ data[095:088] ^ data[103:096] ^
                        data[111:104] ^ data[119:112] ^ data[127:120];
    end
endfunction


// -----------------------------------------------------------------------------
function automatic [7:0] galois_lookup_016;
/*

*/
    input   [7:0]   byte;

    begin case (byte)
        8'h00: galois_lookup_016 = 8'h00;
        8'h01: galois_lookup_016 = 8'h10;
        8'h02: galois_lookup_016 = 8'h20;
        8'h03: galois_lookup_016 = 8'h30;
        8'h04: galois_lookup_016 = 8'h40;
        8'h05: galois_lookup_016 = 8'h50;
        8'h06: galois_lookup_016 = 8'h60;
        8'h07: galois_lookup_016 = 8'h70;
        8'h08: galois_lookup_016 = 8'h80;
        8'h09: galois_lookup_016 = 8'h90;
        8'h0A: galois_lookup_016 = 8'hA0;
        8'h0B: galois_lookup_016 = 8'hB0;
        8'h0C: galois_lookup_016 = 8'hC0;
        8'h0D: galois_lookup_016 = 8'hD0;
        8'h0E: galois_lookup_016 = 8'hE0;
        8'h0F: galois_lookup_016 = 8'hF0;
        8'h10: galois_lookup_016 = 8'hC3;
        8'h11: galois_lookup_016 = 8'hD3;
        8'h12: galois_lookup_016 = 8'hE3;
        8'h13: galois_lookup_016 = 8'hF3;
        8'h14: galois_lookup_016 = 8'h83;
        8'h15: galois_lookup_016 = 8'h93;
        8'h16: galois_lookup_016 = 8'hA3;
        8'h17: galois_lookup_016 = 8'hB3;
        8'h18: galois_lookup_016 = 8'h43;
        8'h19: galois_lookup_016 = 8'h53;
        8'h1A: galois_lookup_016 = 8'h63;
        8'h1B: galois_lookup_016 = 8'h73;
        8'h1C: galois_lookup_016 = 8'h03;
        8'h1D: galois_lookup_016 = 8'h13;
        8'h1E: galois_lookup_016 = 8'h23;
        8'h1F: galois_lookup_016 = 8'h33;
        8'h20: galois_lookup_016 = 8'h45;
        8'h21: galois_lookup_016 = 8'h55;
        8'h22: galois_lookup_016 = 8'h65;
        8'h23: galois_lookup_016 = 8'h75;
        8'h24: galois_lookup_016 = 8'h05;
        8'h25: galois_lookup_016 = 8'h15;
        8'h26: galois_lookup_016 = 8'h25;
        8'h27: galois_lookup_016 = 8'h35;
        8'h28: galois_lookup_016 = 8'hC5;
        8'h29: galois_lookup_016 = 8'hD5;
        8'h2A: galois_lookup_016 = 8'hE5;
        8'h2B: galois_lookup_016 = 8'hF5;
        8'h2C: galois_lookup_016 = 8'h85;
        8'h2D: galois_lookup_016 = 8'h95;
        8'h2E: galois_lookup_016 = 8'hA5;
        8'h2F: galois_lookup_016 = 8'hB5;
        8'h30: galois_lookup_016 = 8'h86;
        8'h31: galois_lookup_016 = 8'h96;
        8'h32: galois_lookup_016 = 8'hA6;
        8'h33: galois_lookup_016 = 8'hB6;
        8'h34: galois_lookup_016 = 8'hC6;
        8'h35: galois_lookup_016 = 8'hD6;
        8'h36: galois_lookup_016 = 8'hE6;
        8'h37: galois_lookup_016 = 8'hF6;
        8'h38: galois_lookup_016 = 8'h06;
        8'h39: galois_lookup_016 = 8'h16;
        8'h3A: galois_lookup_016 = 8'h26;
        8'h3B: galois_lookup_016 = 8'h36;
        8'h3C: galois_lookup_016 = 8'h46;
        8'h3D: galois_lookup_016 = 8'h56;
        8'h3E: galois_lookup_016 = 8'h66;
        8'h3F: galois_lookup_016 = 8'h76;
        8'h40: galois_lookup_016 = 8'h8A;
        8'h41: galois_lookup_016 = 8'h9A;
        8'h42: galois_lookup_016 = 8'hAA;
        8'h43: galois_lookup_016 = 8'hBA;
        8'h44: galois_lookup_016 = 8'hCA;
        8'h45: galois_lookup_016 = 8'hDA;
        8'h46: galois_lookup_016 = 8'hEA;
        8'h47: galois_lookup_016 = 8'hFA;
        8'h48: galois_lookup_016 = 8'h0A;
        8'h49: galois_lookup_016 = 8'h1A;
        8'h4A: galois_lookup_016 = 8'h2A;
        8'h4B: galois_lookup_016 = 8'h3A;
        8'h4C: galois_lookup_016 = 8'h4A;
        8'h4D: galois_lookup_016 = 8'h5A;
        8'h4E: galois_lookup_016 = 8'h6A;
        8'h4F: galois_lookup_016 = 8'h7A;
        8'h50: galois_lookup_016 = 8'h49;
        8'h51: galois_lookup_016 = 8'h59;
        8'h52: galois_lookup_016 = 8'h69;
        8'h53: galois_lookup_016 = 8'h79;
        8'h54: galois_lookup_016 = 8'h09;
        8'h55: galois_lookup_016 = 8'h19;
        8'h56: galois_lookup_016 = 8'h29;
        8'h57: galois_lookup_016 = 8'h39;
        8'h58: galois_lookup_016 = 8'hC9;
        8'h59: galois_lookup_016 = 8'hD9;
        8'h5A: galois_lookup_016 = 8'hE9;
        8'h5B: galois_lookup_016 = 8'hF9;
        8'h5C: galois_lookup_016 = 8'h89;
        8'h5D: galois_lookup_016 = 8'h99;
        8'h5E: galois_lookup_016 = 8'hA9;
        8'h5F: galois_lookup_016 = 8'hB9;
        8'h60: galois_lookup_016 = 8'hCF;
        8'h61: galois_lookup_016 = 8'hDF;
        8'h62: galois_lookup_016 = 8'hEF;
        8'h63: galois_lookup_016 = 8'hFF;
        8'h64: galois_lookup_016 = 8'h8F;
        8'h65: galois_lookup_016 = 8'h9F;
        8'h66: galois_lookup_016 = 8'hAF;
        8'h67: galois_lookup_016 = 8'hBF;
        8'h68: galois_lookup_016 = 8'h4F;
        8'h69: galois_lookup_016 = 8'h5F;
        8'h6A: galois_lookup_016 = 8'h6F;
        8'h6B: galois_lookup_016 = 8'h7F;
        8'h6C: galois_lookup_016 = 8'h0F;
        8'h6D: galois_lookup_016 = 8'h1F;
        8'h6E: galois_lookup_016 = 8'h2F;
        8'h6F: galois_lookup_016 = 8'h3F;
        8'h70: galois_lookup_016 = 8'h0C;
        8'h71: galois_lookup_016 = 8'h1C;
        8'h72: galois_lookup_016 = 8'h2C;
        8'h73: galois_lookup_016 = 8'h3C;
        8'h74: galois_lookup_016 = 8'h4C;
        8'h75: galois_lookup_016 = 8'h5C;
        8'h76: galois_lookup_016 = 8'h6C;
        8'h77: galois_lookup_016 = 8'h7C;
        8'h78: galois_lookup_016 = 8'h8C;
        8'h79: galois_lookup_016 = 8'h9C;
        8'h7A: galois_lookup_016 = 8'hAC;
        8'h7B: galois_lookup_016 = 8'hBC;
        8'h7C: galois_lookup_016 = 8'hCC;
        8'h7D: galois_lookup_016 = 8'hDC;
        8'h7E: galois_lookup_016 = 8'hEC;
        8'h7F: galois_lookup_016 = 8'hFC;
        8'h80: galois_lookup_016 = 8'hD7;
        8'h81: galois_lookup_016 = 8'hC7;
        8'h82: galois_lookup_016 = 8'hF7;
        8'h83: galois_lookup_016 = 8'hE7;
        8'h84: galois_lookup_016 = 8'h97;
        8'h85: galois_lookup_016 = 8'h87;
        8'h86: galois_lookup_016 = 8'hB7;
        8'h87: galois_lookup_016 = 8'hA7;
        8'h88: galois_lookup_016 = 8'h57;
        8'h89: galois_lookup_016 = 8'h47;
        8'h8A: galois_lookup_016 = 8'h77;
        8'h8B: galois_lookup_016 = 8'h67;
        8'h8C: galois_lookup_016 = 8'h17;
        8'h8D: galois_lookup_016 = 8'h07;
        8'h8E: galois_lookup_016 = 8'h37;
        8'h8F: galois_lookup_016 = 8'h27;
        8'h90: galois_lookup_016 = 8'h14;
        8'h91: galois_lookup_016 = 8'h04;
        8'h92: galois_lookup_016 = 8'h34;
        8'h93: galois_lookup_016 = 8'h24;
        8'h94: galois_lookup_016 = 8'h54;
        8'h95: galois_lookup_016 = 8'h44;
        8'h96: galois_lookup_016 = 8'h74;
        8'h97: galois_lookup_016 = 8'h64;
        8'h98: galois_lookup_016 = 8'h94;
        8'h99: galois_lookup_016 = 8'h84;
        8'h9A: galois_lookup_016 = 8'hB4;
        8'h9B: galois_lookup_016 = 8'hA4;
        8'h9C: galois_lookup_016 = 8'hD4;
        8'h9D: galois_lookup_016 = 8'hC4;
        8'h9E: galois_lookup_016 = 8'hF4;
        8'h9F: galois_lookup_016 = 8'hE4;
        8'hA0: galois_lookup_016 = 8'h92;
        8'hA1: galois_lookup_016 = 8'h82;
        8'hA2: galois_lookup_016 = 8'hB2;
        8'hA3: galois_lookup_016 = 8'hA2;
        8'hA4: galois_lookup_016 = 8'hD2;
        8'hA5: galois_lookup_016 = 8'hC2;
        8'hA6: galois_lookup_016 = 8'hF2;
        8'hA7: galois_lookup_016 = 8'hE2;
        8'hA8: galois_lookup_016 = 8'h12;
        8'hA9: galois_lookup_016 = 8'h02;
        8'hAA: galois_lookup_016 = 8'h32;
        8'hAB: galois_lookup_016 = 8'h22;
        8'hAC: galois_lookup_016 = 8'h52;
        8'hAD: galois_lookup_016 = 8'h42;
        8'hAE: galois_lookup_016 = 8'h72;
        8'hAF: galois_lookup_016 = 8'h62;
        8'hB0: galois_lookup_016 = 8'h51;
        8'hB1: galois_lookup_016 = 8'h41;
        8'hB2: galois_lookup_016 = 8'h71;
        8'hB3: galois_lookup_016 = 8'h61;
        8'hB4: galois_lookup_016 = 8'h11;
        8'hB5: galois_lookup_016 = 8'h01;
        8'hB6: galois_lookup_016 = 8'h31;
        8'hB7: galois_lookup_016 = 8'h21;
        8'hB8: galois_lookup_016 = 8'hD1;
        8'hB9: galois_lookup_016 = 8'hC1;
        8'hBA: galois_lookup_016 = 8'hF1;
        8'hBB: galois_lookup_016 = 8'hE1;
        8'hBC: galois_lookup_016 = 8'h91;
        8'hBD: galois_lookup_016 = 8'h81;
        8'hBE: galois_lookup_016 = 8'hB1;
        8'hBF: galois_lookup_016 = 8'hA1;
        8'hC0: galois_lookup_016 = 8'h5D;
        8'hC1: galois_lookup_016 = 8'h4D;
        8'hC2: galois_lookup_016 = 8'h7D;
        8'hC3: galois_lookup_016 = 8'h6D;
        8'hC4: galois_lookup_016 = 8'h1D;
        8'hC5: galois_lookup_016 = 8'h0D;
        8'hC6: galois_lookup_016 = 8'h3D;
        8'hC7: galois_lookup_016 = 8'h2D;
        8'hC8: galois_lookup_016 = 8'hDD;
        8'hC9: galois_lookup_016 = 8'hCD;
        8'hCA: galois_lookup_016 = 8'hFD;
        8'hCB: galois_lookup_016 = 8'hED;
        8'hCC: galois_lookup_016 = 8'h9D;
        8'hCD: galois_lookup_016 = 8'h8D;
        8'hCE: galois_lookup_016 = 8'hBD;
        8'hCF: galois_lookup_016 = 8'hAD;
        8'hD0: galois_lookup_016 = 8'h9E;
        8'hD1: galois_lookup_016 = 8'h8E;
        8'hD2: galois_lookup_016 = 8'hBE;
        8'hD3: galois_lookup_016 = 8'hAE;
        8'hD4: galois_lookup_016 = 8'hDE;
        8'hD5: galois_lookup_016 = 8'hCE;
        8'hD6: galois_lookup_016 = 8'hFE;
        8'hD7: galois_lookup_016 = 8'hEE;
        8'hD8: galois_lookup_016 = 8'h1E;
        8'hD9: galois_lookup_016 = 8'h0E;
        8'hDA: galois_lookup_016 = 8'h3E;
        8'hDB: galois_lookup_016 = 8'h2E;
        8'hDC: galois_lookup_016 = 8'h5E;
        8'hDD: galois_lookup_016 = 8'h4E;
        8'hDE: galois_lookup_016 = 8'h7E;
        8'hDF: galois_lookup_016 = 8'h6E;
        8'hE0: galois_lookup_016 = 8'h18;
        8'hE1: galois_lookup_016 = 8'h08;
        8'hE2: galois_lookup_016 = 8'h38;
        8'hE3: galois_lookup_016 = 8'h28;
        8'hE4: galois_lookup_016 = 8'h58;
        8'hE5: galois_lookup_016 = 8'h48;
        8'hE6: galois_lookup_016 = 8'h78;
        8'hE7: galois_lookup_016 = 8'h68;
        8'hE8: galois_lookup_016 = 8'h98;
        8'hE9: galois_lookup_016 = 8'h88;
        8'hEA: galois_lookup_016 = 8'hB8;
        8'hEB: galois_lookup_016 = 8'hA8;
        8'hEC: galois_lookup_016 = 8'hD8;
        8'hED: galois_lookup_016 = 8'hC8;
        8'hEE: galois_lookup_016 = 8'hF8;
        8'hEF: galois_lookup_016 = 8'hE8;
        8'hF0: galois_lookup_016 = 8'hDB;
        8'hF1: galois_lookup_016 = 8'hCB;
        8'hF2: galois_lookup_016 = 8'hFB;
        8'hF3: galois_lookup_016 = 8'hEB;
        8'hF4: galois_lookup_016 = 8'h9B;
        8'hF5: galois_lookup_016 = 8'h8B;
        8'hF6: galois_lookup_016 = 8'hBB;
        8'hF7: galois_lookup_016 = 8'hAB;
        8'hF8: galois_lookup_016 = 8'h5B;
        8'hF9: galois_lookup_016 = 8'h4B;
        8'hFA: galois_lookup_016 = 8'h7B;
        8'hFB: galois_lookup_016 = 8'h6B;
        8'hFC: galois_lookup_016 = 8'h1B;
        8'hFD: galois_lookup_016 = 8'h0B;
        8'hFE: galois_lookup_016 = 8'h3B;
        8'hFF: galois_lookup_016 = 8'h2B;
    endcase end
endfunction

// -----------------------------------------------------------------------------
function automatic [7:0] galois_lookup_032;
/*

*/
    input   [7:0]   byte;

    begin case (byte)
        8'h00: galois_lookup_032 = 8'h00;
        8'h01: galois_lookup_032 = 8'h20;
        8'h02: galois_lookup_032 = 8'h40;
        8'h03: galois_lookup_032 = 8'h60;
        8'h04: galois_lookup_032 = 8'h80;
        8'h05: galois_lookup_032 = 8'hA0;
        8'h06: galois_lookup_032 = 8'hC0;
        8'h07: galois_lookup_032 = 8'hE0;
        8'h08: galois_lookup_032 = 8'hC3;
        8'h09: galois_lookup_032 = 8'hE3;
        8'h0A: galois_lookup_032 = 8'h83;
        8'h0B: galois_lookup_032 = 8'hA3;
        8'h0C: galois_lookup_032 = 8'h43;
        8'h0D: galois_lookup_032 = 8'h63;
        8'h0E: galois_lookup_032 = 8'h03;
        8'h0F: galois_lookup_032 = 8'h23;
        8'h10: galois_lookup_032 = 8'h45;
        8'h11: galois_lookup_032 = 8'h65;
        8'h12: galois_lookup_032 = 8'h05;
        8'h13: galois_lookup_032 = 8'h25;
        8'h14: galois_lookup_032 = 8'hC5;
        8'h15: galois_lookup_032 = 8'hE5;
        8'h16: galois_lookup_032 = 8'h85;
        8'h17: galois_lookup_032 = 8'hA5;
        8'h18: galois_lookup_032 = 8'h86;
        8'h19: galois_lookup_032 = 8'hA6;
        8'h1A: galois_lookup_032 = 8'hC6;
        8'h1B: galois_lookup_032 = 8'hE6;
        8'h1C: galois_lookup_032 = 8'h06;
        8'h1D: galois_lookup_032 = 8'h26;
        8'h1E: galois_lookup_032 = 8'h46;
        8'h1F: galois_lookup_032 = 8'h66;
        8'h20: galois_lookup_032 = 8'h8A;
        8'h21: galois_lookup_032 = 8'hAA;
        8'h22: galois_lookup_032 = 8'hCA;
        8'h23: galois_lookup_032 = 8'hEA;
        8'h24: galois_lookup_032 = 8'h0A;
        8'h25: galois_lookup_032 = 8'h2A;
        8'h26: galois_lookup_032 = 8'h4A;
        8'h27: galois_lookup_032 = 8'h6A;
        8'h28: galois_lookup_032 = 8'h49;
        8'h29: galois_lookup_032 = 8'h69;
        8'h2A: galois_lookup_032 = 8'h09;
        8'h2B: galois_lookup_032 = 8'h29;
        8'h2C: galois_lookup_032 = 8'hC9;
        8'h2D: galois_lookup_032 = 8'hE9;
        8'h2E: galois_lookup_032 = 8'h89;
        8'h2F: galois_lookup_032 = 8'hA9;
        8'h30: galois_lookup_032 = 8'hCF;
        8'h31: galois_lookup_032 = 8'hEF;
        8'h32: galois_lookup_032 = 8'h8F;
        8'h33: galois_lookup_032 = 8'hAF;
        8'h34: galois_lookup_032 = 8'h4F;
        8'h35: galois_lookup_032 = 8'h6F;
        8'h36: galois_lookup_032 = 8'h0F;
        8'h37: galois_lookup_032 = 8'h2F;
        8'h38: galois_lookup_032 = 8'h0C;
        8'h39: galois_lookup_032 = 8'h2C;
        8'h3A: galois_lookup_032 = 8'h4C;
        8'h3B: galois_lookup_032 = 8'h6C;
        8'h3C: galois_lookup_032 = 8'h8C;
        8'h3D: galois_lookup_032 = 8'hAC;
        8'h3E: galois_lookup_032 = 8'hCC;
        8'h3F: galois_lookup_032 = 8'hEC;
        8'h40: galois_lookup_032 = 8'hD7;
        8'h41: galois_lookup_032 = 8'hF7;
        8'h42: galois_lookup_032 = 8'h97;
        8'h43: galois_lookup_032 = 8'hB7;
        8'h44: galois_lookup_032 = 8'h57;
        8'h45: galois_lookup_032 = 8'h77;
        8'h46: galois_lookup_032 = 8'h17;
        8'h47: galois_lookup_032 = 8'h37;
        8'h48: galois_lookup_032 = 8'h14;
        8'h49: galois_lookup_032 = 8'h34;
        8'h4A: galois_lookup_032 = 8'h54;
        8'h4B: galois_lookup_032 = 8'h74;
        8'h4C: galois_lookup_032 = 8'h94;
        8'h4D: galois_lookup_032 = 8'hB4;
        8'h4E: galois_lookup_032 = 8'hD4;
        8'h4F: galois_lookup_032 = 8'hF4;
        8'h50: galois_lookup_032 = 8'h92;
        8'h51: galois_lookup_032 = 8'hB2;
        8'h52: galois_lookup_032 = 8'hD2;
        8'h53: galois_lookup_032 = 8'hF2;
        8'h54: galois_lookup_032 = 8'h12;
        8'h55: galois_lookup_032 = 8'h32;
        8'h56: galois_lookup_032 = 8'h52;
        8'h57: galois_lookup_032 = 8'h72;
        8'h58: galois_lookup_032 = 8'h51;
        8'h59: galois_lookup_032 = 8'h71;
        8'h5A: galois_lookup_032 = 8'h11;
        8'h5B: galois_lookup_032 = 8'h31;
        8'h5C: galois_lookup_032 = 8'hD1;
        8'h5D: galois_lookup_032 = 8'hF1;
        8'h5E: galois_lookup_032 = 8'h91;
        8'h5F: galois_lookup_032 = 8'hB1;
        8'h60: galois_lookup_032 = 8'h5D;
        8'h61: galois_lookup_032 = 8'h7D;
        8'h62: galois_lookup_032 = 8'h1D;
        8'h63: galois_lookup_032 = 8'h3D;
        8'h64: galois_lookup_032 = 8'hDD;
        8'h65: galois_lookup_032 = 8'hFD;
        8'h66: galois_lookup_032 = 8'h9D;
        8'h67: galois_lookup_032 = 8'hBD;
        8'h68: galois_lookup_032 = 8'h9E;
        8'h69: galois_lookup_032 = 8'hBE;
        8'h6A: galois_lookup_032 = 8'hDE;
        8'h6B: galois_lookup_032 = 8'hFE;
        8'h6C: galois_lookup_032 = 8'h1E;
        8'h6D: galois_lookup_032 = 8'h3E;
        8'h6E: galois_lookup_032 = 8'h5E;
        8'h6F: galois_lookup_032 = 8'h7E;
        8'h70: galois_lookup_032 = 8'h18;
        8'h71: galois_lookup_032 = 8'h38;
        8'h72: galois_lookup_032 = 8'h58;
        8'h73: galois_lookup_032 = 8'h78;
        8'h74: galois_lookup_032 = 8'h98;
        8'h75: galois_lookup_032 = 8'hB8;
        8'h76: galois_lookup_032 = 8'hD8;
        8'h77: galois_lookup_032 = 8'hF8;
        8'h78: galois_lookup_032 = 8'hDB;
        8'h79: galois_lookup_032 = 8'hFB;
        8'h7A: galois_lookup_032 = 8'h9B;
        8'h7B: galois_lookup_032 = 8'hBB;
        8'h7C: galois_lookup_032 = 8'h5B;
        8'h7D: galois_lookup_032 = 8'h7B;
        8'h7E: galois_lookup_032 = 8'h1B;
        8'h7F: galois_lookup_032 = 8'h3B;
        8'h80: galois_lookup_032 = 8'h6D;
        8'h81: galois_lookup_032 = 8'h4D;
        8'h82: galois_lookup_032 = 8'h2D;
        8'h83: galois_lookup_032 = 8'h0D;
        8'h84: galois_lookup_032 = 8'hED;
        8'h85: galois_lookup_032 = 8'hCD;
        8'h86: galois_lookup_032 = 8'hAD;
        8'h87: galois_lookup_032 = 8'h8D;
        8'h88: galois_lookup_032 = 8'hAE;
        8'h89: galois_lookup_032 = 8'h8E;
        8'h8A: galois_lookup_032 = 8'hEE;
        8'h8B: galois_lookup_032 = 8'hCE;
        8'h8C: galois_lookup_032 = 8'h2E;
        8'h8D: galois_lookup_032 = 8'h0E;
        8'h8E: galois_lookup_032 = 8'h6E;
        8'h8F: galois_lookup_032 = 8'h4E;
        8'h90: galois_lookup_032 = 8'h28;
        8'h91: galois_lookup_032 = 8'h08;
        8'h92: galois_lookup_032 = 8'h68;
        8'h93: galois_lookup_032 = 8'h48;
        8'h94: galois_lookup_032 = 8'hA8;
        8'h95: galois_lookup_032 = 8'h88;
        8'h96: galois_lookup_032 = 8'hE8;
        8'h97: galois_lookup_032 = 8'hC8;
        8'h98: galois_lookup_032 = 8'hEB;
        8'h99: galois_lookup_032 = 8'hCB;
        8'h9A: galois_lookup_032 = 8'hAB;
        8'h9B: galois_lookup_032 = 8'h8B;
        8'h9C: galois_lookup_032 = 8'h6B;
        8'h9D: galois_lookup_032 = 8'h4B;
        8'h9E: galois_lookup_032 = 8'h2B;
        8'h9F: galois_lookup_032 = 8'h0B;
        8'hA0: galois_lookup_032 = 8'hE7;
        8'hA1: galois_lookup_032 = 8'hC7;
        8'hA2: galois_lookup_032 = 8'hA7;
        8'hA3: galois_lookup_032 = 8'h87;
        8'hA4: galois_lookup_032 = 8'h67;
        8'hA5: galois_lookup_032 = 8'h47;
        8'hA6: galois_lookup_032 = 8'h27;
        8'hA7: galois_lookup_032 = 8'h07;
        8'hA8: galois_lookup_032 = 8'h24;
        8'hA9: galois_lookup_032 = 8'h04;
        8'hAA: galois_lookup_032 = 8'h64;
        8'hAB: galois_lookup_032 = 8'h44;
        8'hAC: galois_lookup_032 = 8'hA4;
        8'hAD: galois_lookup_032 = 8'h84;
        8'hAE: galois_lookup_032 = 8'hE4;
        8'hAF: galois_lookup_032 = 8'hC4;
        8'hB0: galois_lookup_032 = 8'hA2;
        8'hB1: galois_lookup_032 = 8'h82;
        8'hB2: galois_lookup_032 = 8'hE2;
        8'hB3: galois_lookup_032 = 8'hC2;
        8'hB4: galois_lookup_032 = 8'h22;
        8'hB5: galois_lookup_032 = 8'h02;
        8'hB6: galois_lookup_032 = 8'h62;
        8'hB7: galois_lookup_032 = 8'h42;
        8'hB8: galois_lookup_032 = 8'h61;
        8'hB9: galois_lookup_032 = 8'h41;
        8'hBA: galois_lookup_032 = 8'h21;
        8'hBB: galois_lookup_032 = 8'h01;
        8'hBC: galois_lookup_032 = 8'hE1;
        8'hBD: galois_lookup_032 = 8'hC1;
        8'hBE: galois_lookup_032 = 8'hA1;
        8'hBF: galois_lookup_032 = 8'h81;
        8'hC0: galois_lookup_032 = 8'hBA;
        8'hC1: galois_lookup_032 = 8'h9A;
        8'hC2: galois_lookup_032 = 8'hFA;
        8'hC3: galois_lookup_032 = 8'hDA;
        8'hC4: galois_lookup_032 = 8'h3A;
        8'hC5: galois_lookup_032 = 8'h1A;
        8'hC6: galois_lookup_032 = 8'h7A;
        8'hC7: galois_lookup_032 = 8'h5A;
        8'hC8: galois_lookup_032 = 8'h79;
        8'hC9: galois_lookup_032 = 8'h59;
        8'hCA: galois_lookup_032 = 8'h39;
        8'hCB: galois_lookup_032 = 8'h19;
        8'hCC: galois_lookup_032 = 8'hF9;
        8'hCD: galois_lookup_032 = 8'hD9;
        8'hCE: galois_lookup_032 = 8'hB9;
        8'hCF: galois_lookup_032 = 8'h99;
        8'hD0: galois_lookup_032 = 8'hFF;
        8'hD1: galois_lookup_032 = 8'hDF;
        8'hD2: galois_lookup_032 = 8'hBF;
        8'hD3: galois_lookup_032 = 8'h9F;
        8'hD4: galois_lookup_032 = 8'h7F;
        8'hD5: galois_lookup_032 = 8'h5F;
        8'hD6: galois_lookup_032 = 8'h3F;
        8'hD7: galois_lookup_032 = 8'h1F;
        8'hD8: galois_lookup_032 = 8'h3C;
        8'hD9: galois_lookup_032 = 8'h1C;
        8'hDA: galois_lookup_032 = 8'h7C;
        8'hDB: galois_lookup_032 = 8'h5C;
        8'hDC: galois_lookup_032 = 8'hBC;
        8'hDD: galois_lookup_032 = 8'h9C;
        8'hDE: galois_lookup_032 = 8'hFC;
        8'hDF: galois_lookup_032 = 8'hDC;
        8'hE0: galois_lookup_032 = 8'h30;
        8'hE1: galois_lookup_032 = 8'h10;
        8'hE2: galois_lookup_032 = 8'h70;
        8'hE3: galois_lookup_032 = 8'h50;
        8'hE4: galois_lookup_032 = 8'hB0;
        8'hE5: galois_lookup_032 = 8'h90;
        8'hE6: galois_lookup_032 = 8'hF0;
        8'hE7: galois_lookup_032 = 8'hD0;
        8'hE8: galois_lookup_032 = 8'hF3;
        8'hE9: galois_lookup_032 = 8'hD3;
        8'hEA: galois_lookup_032 = 8'hB3;
        8'hEB: galois_lookup_032 = 8'h93;
        8'hEC: galois_lookup_032 = 8'h73;
        8'hED: galois_lookup_032 = 8'h53;
        8'hEE: galois_lookup_032 = 8'h33;
        8'hEF: galois_lookup_032 = 8'h13;
        8'hF0: galois_lookup_032 = 8'h75;
        8'hF1: galois_lookup_032 = 8'h55;
        8'hF2: galois_lookup_032 = 8'h35;
        8'hF3: galois_lookup_032 = 8'h15;
        8'hF4: galois_lookup_032 = 8'hF5;
        8'hF5: galois_lookup_032 = 8'hD5;
        8'hF6: galois_lookup_032 = 8'hB5;
        8'hF7: galois_lookup_032 = 8'h95;
        8'hF8: galois_lookup_032 = 8'hB6;
        8'hF9: galois_lookup_032 = 8'h96;
        8'hFA: galois_lookup_032 = 8'hF6;
        8'hFB: galois_lookup_032 = 8'hD6;
        8'hFC: galois_lookup_032 = 8'h36;
        8'hFD: galois_lookup_032 = 8'h16;
        8'hFE: galois_lookup_032 = 8'h76;
        8'hFF: galois_lookup_032 = 8'h56;
    endcase end
endfunction

// -----------------------------------------------------------------------------
function automatic [7:0] galois_lookup_133;
/*

*/
    input   [7:0]   byte;

    begin case (byte)
        8'h00: galois_lookup_133 = 8'h00;
        8'h01: galois_lookup_133 = 8'h85;
        8'h02: galois_lookup_133 = 8'hC9;
        8'h03: galois_lookup_133 = 8'h4C;
        8'h04: galois_lookup_133 = 8'h51;
        8'h05: galois_lookup_133 = 8'hD4;
        8'h06: galois_lookup_133 = 8'h98;
        8'h07: galois_lookup_133 = 8'h1D;
        8'h08: galois_lookup_133 = 8'hA2;
        8'h09: galois_lookup_133 = 8'h27;
        8'h0A: galois_lookup_133 = 8'h6B;
        8'h0B: galois_lookup_133 = 8'hEE;
        8'h0C: galois_lookup_133 = 8'hF3;
        8'h0D: galois_lookup_133 = 8'h76;
        8'h0E: galois_lookup_133 = 8'h3A;
        8'h0F: galois_lookup_133 = 8'hBF;
        8'h10: galois_lookup_133 = 8'h87;
        8'h11: galois_lookup_133 = 8'h02;
        8'h12: galois_lookup_133 = 8'h4E;
        8'h13: galois_lookup_133 = 8'hCB;
        8'h14: galois_lookup_133 = 8'hD6;
        8'h15: galois_lookup_133 = 8'h53;
        8'h16: galois_lookup_133 = 8'h1F;
        8'h17: galois_lookup_133 = 8'h9A;
        8'h18: galois_lookup_133 = 8'h25;
        8'h19: galois_lookup_133 = 8'hA0;
        8'h1A: galois_lookup_133 = 8'hEC;
        8'h1B: galois_lookup_133 = 8'h69;
        8'h1C: galois_lookup_133 = 8'h74;
        8'h1D: galois_lookup_133 = 8'hF1;
        8'h1E: galois_lookup_133 = 8'hBD;
        8'h1F: galois_lookup_133 = 8'h38;
        8'h20: galois_lookup_133 = 8'hCD;
        8'h21: galois_lookup_133 = 8'h48;
        8'h22: galois_lookup_133 = 8'h04;
        8'h23: galois_lookup_133 = 8'h81;
        8'h24: galois_lookup_133 = 8'h9C;
        8'h25: galois_lookup_133 = 8'h19;
        8'h26: galois_lookup_133 = 8'h55;
        8'h27: galois_lookup_133 = 8'hD0;
        8'h28: galois_lookup_133 = 8'h6F;
        8'h29: galois_lookup_133 = 8'hEA;
        8'h2A: galois_lookup_133 = 8'hA6;
        8'h2B: galois_lookup_133 = 8'h23;
        8'h2C: galois_lookup_133 = 8'h3E;
        8'h2D: galois_lookup_133 = 8'hBB;
        8'h2E: galois_lookup_133 = 8'hF7;
        8'h2F: galois_lookup_133 = 8'h72;
        8'h30: galois_lookup_133 = 8'h4A;
        8'h31: galois_lookup_133 = 8'hCF;
        8'h32: galois_lookup_133 = 8'h83;
        8'h33: galois_lookup_133 = 8'h06;
        8'h34: galois_lookup_133 = 8'h1B;
        8'h35: galois_lookup_133 = 8'h9E;
        8'h36: galois_lookup_133 = 8'hD2;
        8'h37: galois_lookup_133 = 8'h57;
        8'h38: galois_lookup_133 = 8'hE8;
        8'h39: galois_lookup_133 = 8'h6D;
        8'h3A: galois_lookup_133 = 8'h21;
        8'h3B: galois_lookup_133 = 8'hA4;
        8'h3C: galois_lookup_133 = 8'hB9;
        8'h3D: galois_lookup_133 = 8'h3C;
        8'h3E: galois_lookup_133 = 8'h70;
        8'h3F: galois_lookup_133 = 8'hF5;
        8'h40: galois_lookup_133 = 8'h59;
        8'h41: galois_lookup_133 = 8'hDC;
        8'h42: galois_lookup_133 = 8'h90;
        8'h43: galois_lookup_133 = 8'h15;
        8'h44: galois_lookup_133 = 8'h08;
        8'h45: galois_lookup_133 = 8'h8D;
        8'h46: galois_lookup_133 = 8'hC1;
        8'h47: galois_lookup_133 = 8'h44;
        8'h48: galois_lookup_133 = 8'hFB;
        8'h49: galois_lookup_133 = 8'h7E;
        8'h4A: galois_lookup_133 = 8'h32;
        8'h4B: galois_lookup_133 = 8'hB7;
        8'h4C: galois_lookup_133 = 8'hAA;
        8'h4D: galois_lookup_133 = 8'h2F;
        8'h4E: galois_lookup_133 = 8'h63;
        8'h4F: galois_lookup_133 = 8'hE6;
        8'h50: galois_lookup_133 = 8'hDE;
        8'h51: galois_lookup_133 = 8'h5B;
        8'h52: galois_lookup_133 = 8'h17;
        8'h53: galois_lookup_133 = 8'h92;
        8'h54: galois_lookup_133 = 8'h8F;
        8'h55: galois_lookup_133 = 8'h0A;
        8'h56: galois_lookup_133 = 8'h46;
        8'h57: galois_lookup_133 = 8'hC3;
        8'h58: galois_lookup_133 = 8'h7C;
        8'h59: galois_lookup_133 = 8'hF9;
        8'h5A: galois_lookup_133 = 8'hB5;
        8'h5B: galois_lookup_133 = 8'h30;
        8'h5C: galois_lookup_133 = 8'h2D;
        8'h5D: galois_lookup_133 = 8'hA8;
        8'h5E: galois_lookup_133 = 8'hE4;
        8'h5F: galois_lookup_133 = 8'h61;
        8'h60: galois_lookup_133 = 8'h94;
        8'h61: galois_lookup_133 = 8'h11;
        8'h62: galois_lookup_133 = 8'h5D;
        8'h63: galois_lookup_133 = 8'hD8;
        8'h64: galois_lookup_133 = 8'hC5;
        8'h65: galois_lookup_133 = 8'h40;
        8'h66: galois_lookup_133 = 8'h0C;
        8'h67: galois_lookup_133 = 8'h89;
        8'h68: galois_lookup_133 = 8'h36;
        8'h69: galois_lookup_133 = 8'hB3;
        8'h6A: galois_lookup_133 = 8'hFF;
        8'h6B: galois_lookup_133 = 8'h7A;
        8'h6C: galois_lookup_133 = 8'h67;
        8'h6D: galois_lookup_133 = 8'hE2;
        8'h6E: galois_lookup_133 = 8'hAE;
        8'h6F: galois_lookup_133 = 8'h2B;
        8'h70: galois_lookup_133 = 8'h13;
        8'h71: galois_lookup_133 = 8'h96;
        8'h72: galois_lookup_133 = 8'hDA;
        8'h73: galois_lookup_133 = 8'h5F;
        8'h74: galois_lookup_133 = 8'h42;
        8'h75: galois_lookup_133 = 8'hC7;
        8'h76: galois_lookup_133 = 8'h8B;
        8'h77: galois_lookup_133 = 8'h0E;
        8'h78: galois_lookup_133 = 8'hB1;
        8'h79: galois_lookup_133 = 8'h34;
        8'h7A: galois_lookup_133 = 8'h78;
        8'h7B: galois_lookup_133 = 8'hFD;
        8'h7C: galois_lookup_133 = 8'hE0;
        8'h7D: galois_lookup_133 = 8'h65;
        8'h7E: galois_lookup_133 = 8'h29;
        8'h7F: galois_lookup_133 = 8'hAC;
        8'h80: galois_lookup_133 = 8'hB2;
        8'h81: galois_lookup_133 = 8'h37;
        8'h82: galois_lookup_133 = 8'h7B;
        8'h83: galois_lookup_133 = 8'hFE;
        8'h84: galois_lookup_133 = 8'hE3;
        8'h85: galois_lookup_133 = 8'h66;
        8'h86: galois_lookup_133 = 8'h2A;
        8'h87: galois_lookup_133 = 8'hAF;
        8'h88: galois_lookup_133 = 8'h10;
        8'h89: galois_lookup_133 = 8'h95;
        8'h8A: galois_lookup_133 = 8'hD9;
        8'h8B: galois_lookup_133 = 8'h5C;
        8'h8C: galois_lookup_133 = 8'h41;
        8'h8D: galois_lookup_133 = 8'hC4;
        8'h8E: galois_lookup_133 = 8'h88;
        8'h8F: galois_lookup_133 = 8'h0D;
        8'h90: galois_lookup_133 = 8'h35;
        8'h91: galois_lookup_133 = 8'hB0;
        8'h92: galois_lookup_133 = 8'hFC;
        8'h93: galois_lookup_133 = 8'h79;
        8'h94: galois_lookup_133 = 8'h64;
        8'h95: galois_lookup_133 = 8'hE1;
        8'h96: galois_lookup_133 = 8'hAD;
        8'h97: galois_lookup_133 = 8'h28;
        8'h98: galois_lookup_133 = 8'h97;
        8'h99: galois_lookup_133 = 8'h12;
        8'h9A: galois_lookup_133 = 8'h5E;
        8'h9B: galois_lookup_133 = 8'hDB;
        8'h9C: galois_lookup_133 = 8'hC6;
        8'h9D: galois_lookup_133 = 8'h43;
        8'h9E: galois_lookup_133 = 8'h0F;
        8'h9F: galois_lookup_133 = 8'h8A;
        8'hA0: galois_lookup_133 = 8'h7F;
        8'hA1: galois_lookup_133 = 8'hFA;
        8'hA2: galois_lookup_133 = 8'hB6;
        8'hA3: galois_lookup_133 = 8'h33;
        8'hA4: galois_lookup_133 = 8'h2E;
        8'hA5: galois_lookup_133 = 8'hAB;
        8'hA6: galois_lookup_133 = 8'hE7;
        8'hA7: galois_lookup_133 = 8'h62;
        8'hA8: galois_lookup_133 = 8'hDD;
        8'hA9: galois_lookup_133 = 8'h58;
        8'hAA: galois_lookup_133 = 8'h14;
        8'hAB: galois_lookup_133 = 8'h91;
        8'hAC: galois_lookup_133 = 8'h8C;
        8'hAD: galois_lookup_133 = 8'h09;
        8'hAE: galois_lookup_133 = 8'h45;
        8'hAF: galois_lookup_133 = 8'hC0;
        8'hB0: galois_lookup_133 = 8'hF8;
        8'hB1: galois_lookup_133 = 8'h7D;
        8'hB2: galois_lookup_133 = 8'h31;
        8'hB3: galois_lookup_133 = 8'hB4;
        8'hB4: galois_lookup_133 = 8'hA9;
        8'hB5: galois_lookup_133 = 8'h2C;
        8'hB6: galois_lookup_133 = 8'h60;
        8'hB7: galois_lookup_133 = 8'hE5;
        8'hB8: galois_lookup_133 = 8'h5A;
        8'hB9: galois_lookup_133 = 8'hDF;
        8'hBA: galois_lookup_133 = 8'h93;
        8'hBB: galois_lookup_133 = 8'h16;
        8'hBC: galois_lookup_133 = 8'h0B;
        8'hBD: galois_lookup_133 = 8'h8E;
        8'hBE: galois_lookup_133 = 8'hC2;
        8'hBF: galois_lookup_133 = 8'h47;
        8'hC0: galois_lookup_133 = 8'hEB;
        8'hC1: galois_lookup_133 = 8'h6E;
        8'hC2: galois_lookup_133 = 8'h22;
        8'hC3: galois_lookup_133 = 8'hA7;
        8'hC4: galois_lookup_133 = 8'hBA;
        8'hC5: galois_lookup_133 = 8'h3F;
        8'hC6: galois_lookup_133 = 8'h73;
        8'hC7: galois_lookup_133 = 8'hF6;
        8'hC8: galois_lookup_133 = 8'h49;
        8'hC9: galois_lookup_133 = 8'hCC;
        8'hCA: galois_lookup_133 = 8'h80;
        8'hCB: galois_lookup_133 = 8'h05;
        8'hCC: galois_lookup_133 = 8'h18;
        8'hCD: galois_lookup_133 = 8'h9D;
        8'hCE: galois_lookup_133 = 8'hD1;
        8'hCF: galois_lookup_133 = 8'h54;
        8'hD0: galois_lookup_133 = 8'h6C;
        8'hD1: galois_lookup_133 = 8'hE9;
        8'hD2: galois_lookup_133 = 8'hA5;
        8'hD3: galois_lookup_133 = 8'h20;
        8'hD4: galois_lookup_133 = 8'h3D;
        8'hD5: galois_lookup_133 = 8'hB8;
        8'hD6: galois_lookup_133 = 8'hF4;
        8'hD7: galois_lookup_133 = 8'h71;
        8'hD8: galois_lookup_133 = 8'hCE;
        8'hD9: galois_lookup_133 = 8'h4B;
        8'hDA: galois_lookup_133 = 8'h07;
        8'hDB: galois_lookup_133 = 8'h82;
        8'hDC: galois_lookup_133 = 8'h9F;
        8'hDD: galois_lookup_133 = 8'h1A;
        8'hDE: galois_lookup_133 = 8'h56;
        8'hDF: galois_lookup_133 = 8'hD3;
        8'hE0: galois_lookup_133 = 8'h26;
        8'hE1: galois_lookup_133 = 8'hA3;
        8'hE2: galois_lookup_133 = 8'hEF;
        8'hE3: galois_lookup_133 = 8'h6A;
        8'hE4: galois_lookup_133 = 8'h77;
        8'hE5: galois_lookup_133 = 8'hF2;
        8'hE6: galois_lookup_133 = 8'hBE;
        8'hE7: galois_lookup_133 = 8'h3B;
        8'hE8: galois_lookup_133 = 8'h84;
        8'hE9: galois_lookup_133 = 8'h01;
        8'hEA: galois_lookup_133 = 8'h4D;
        8'hEB: galois_lookup_133 = 8'hC8;
        8'hEC: galois_lookup_133 = 8'hD5;
        8'hED: galois_lookup_133 = 8'h50;
        8'hEE: galois_lookup_133 = 8'h1C;
        8'hEF: galois_lookup_133 = 8'h99;
        8'hF0: galois_lookup_133 = 8'hA1;
        8'hF1: galois_lookup_133 = 8'h24;
        8'hF2: galois_lookup_133 = 8'h68;
        8'hF3: galois_lookup_133 = 8'hED;
        8'hF4: galois_lookup_133 = 8'hF0;
        8'hF5: galois_lookup_133 = 8'h75;
        8'hF6: galois_lookup_133 = 8'h39;
        8'hF7: galois_lookup_133 = 8'hBC;
        8'hF8: galois_lookup_133 = 8'h03;
        8'hF9: galois_lookup_133 = 8'h86;
        8'hFA: galois_lookup_133 = 8'hCA;
        8'hFB: galois_lookup_133 = 8'h4F;
        8'hFC: galois_lookup_133 = 8'h52;
        8'hFD: galois_lookup_133 = 8'hD7;
        8'hFE: galois_lookup_133 = 8'h9B;
        8'hFF: galois_lookup_133 = 8'h1E;
    endcase end
endfunction

// -----------------------------------------------------------------------------
function automatic [7:0] galois_lookup_148;
/*

*/
    input   [7:0]   byte;

    begin case (byte)
        8'h00: galois_lookup_148 = 8'h00;
        8'h01: galois_lookup_148 = 8'h94;
        8'h02: galois_lookup_148 = 8'hEB;
        8'h03: galois_lookup_148 = 8'h7F;
        8'h04: galois_lookup_148 = 8'h15;
        8'h05: galois_lookup_148 = 8'h81;
        8'h06: galois_lookup_148 = 8'hFE;
        8'h07: galois_lookup_148 = 8'h6A;
        8'h08: galois_lookup_148 = 8'h2A;
        8'h09: galois_lookup_148 = 8'hBE;
        8'h0A: galois_lookup_148 = 8'hC1;
        8'h0B: galois_lookup_148 = 8'h55;
        8'h0C: galois_lookup_148 = 8'h3F;
        8'h0D: galois_lookup_148 = 8'hAB;
        8'h0E: galois_lookup_148 = 8'hD4;
        8'h0F: galois_lookup_148 = 8'h40;
        8'h10: galois_lookup_148 = 8'h54;
        8'h11: galois_lookup_148 = 8'hC0;
        8'h12: galois_lookup_148 = 8'hBF;
        8'h13: galois_lookup_148 = 8'h2B;
        8'h14: galois_lookup_148 = 8'h41;
        8'h15: galois_lookup_148 = 8'hD5;
        8'h16: galois_lookup_148 = 8'hAA;
        8'h17: galois_lookup_148 = 8'h3E;
        8'h18: galois_lookup_148 = 8'h7E;
        8'h19: galois_lookup_148 = 8'hEA;
        8'h1A: galois_lookup_148 = 8'h95;
        8'h1B: galois_lookup_148 = 8'h01;
        8'h1C: galois_lookup_148 = 8'h6B;
        8'h1D: galois_lookup_148 = 8'hFF;
        8'h1E: galois_lookup_148 = 8'h80;
        8'h1F: galois_lookup_148 = 8'h14;
        8'h20: galois_lookup_148 = 8'hA8;
        8'h21: galois_lookup_148 = 8'h3C;
        8'h22: galois_lookup_148 = 8'h43;
        8'h23: galois_lookup_148 = 8'hD7;
        8'h24: galois_lookup_148 = 8'hBD;
        8'h25: galois_lookup_148 = 8'h29;
        8'h26: galois_lookup_148 = 8'h56;
        8'h27: galois_lookup_148 = 8'hC2;
        8'h28: galois_lookup_148 = 8'h82;
        8'h29: galois_lookup_148 = 8'h16;
        8'h2A: galois_lookup_148 = 8'h69;
        8'h2B: galois_lookup_148 = 8'hFD;
        8'h2C: galois_lookup_148 = 8'h97;
        8'h2D: galois_lookup_148 = 8'h03;
        8'h2E: galois_lookup_148 = 8'h7C;
        8'h2F: galois_lookup_148 = 8'hE8;
        8'h30: galois_lookup_148 = 8'hFC;
        8'h31: galois_lookup_148 = 8'h68;
        8'h32: galois_lookup_148 = 8'h17;
        8'h33: galois_lookup_148 = 8'h83;
        8'h34: galois_lookup_148 = 8'hE9;
        8'h35: galois_lookup_148 = 8'h7D;
        8'h36: galois_lookup_148 = 8'h02;
        8'h37: galois_lookup_148 = 8'h96;
        8'h38: galois_lookup_148 = 8'hD6;
        8'h39: galois_lookup_148 = 8'h42;
        8'h3A: galois_lookup_148 = 8'h3D;
        8'h3B: galois_lookup_148 = 8'hA9;
        8'h3C: galois_lookup_148 = 8'hC3;
        8'h3D: galois_lookup_148 = 8'h57;
        8'h3E: galois_lookup_148 = 8'h28;
        8'h3F: galois_lookup_148 = 8'hBC;
        8'h40: galois_lookup_148 = 8'h93;
        8'h41: galois_lookup_148 = 8'h07;
        8'h42: galois_lookup_148 = 8'h78;
        8'h43: galois_lookup_148 = 8'hEC;
        8'h44: galois_lookup_148 = 8'h86;
        8'h45: galois_lookup_148 = 8'h12;
        8'h46: galois_lookup_148 = 8'h6D;
        8'h47: galois_lookup_148 = 8'hF9;
        8'h48: galois_lookup_148 = 8'hB9;
        8'h49: galois_lookup_148 = 8'h2D;
        8'h4A: galois_lookup_148 = 8'h52;
        8'h4B: galois_lookup_148 = 8'hC6;
        8'h4C: galois_lookup_148 = 8'hAC;
        8'h4D: galois_lookup_148 = 8'h38;
        8'h4E: galois_lookup_148 = 8'h47;
        8'h4F: galois_lookup_148 = 8'hD3;
        8'h50: galois_lookup_148 = 8'hC7;
        8'h51: galois_lookup_148 = 8'h53;
        8'h52: galois_lookup_148 = 8'h2C;
        8'h53: galois_lookup_148 = 8'hB8;
        8'h54: galois_lookup_148 = 8'hD2;
        8'h55: galois_lookup_148 = 8'h46;
        8'h56: galois_lookup_148 = 8'h39;
        8'h57: galois_lookup_148 = 8'hAD;
        8'h58: galois_lookup_148 = 8'hED;
        8'h59: galois_lookup_148 = 8'h79;
        8'h5A: galois_lookup_148 = 8'h06;
        8'h5B: galois_lookup_148 = 8'h92;
        8'h5C: galois_lookup_148 = 8'hF8;
        8'h5D: galois_lookup_148 = 8'h6C;
        8'h5E: galois_lookup_148 = 8'h13;
        8'h5F: galois_lookup_148 = 8'h87;
        8'h60: galois_lookup_148 = 8'h3B;
        8'h61: galois_lookup_148 = 8'hAF;
        8'h62: galois_lookup_148 = 8'hD0;
        8'h63: galois_lookup_148 = 8'h44;
        8'h64: galois_lookup_148 = 8'h2E;
        8'h65: galois_lookup_148 = 8'hBA;
        8'h66: galois_lookup_148 = 8'hC5;
        8'h67: galois_lookup_148 = 8'h51;
        8'h68: galois_lookup_148 = 8'h11;
        8'h69: galois_lookup_148 = 8'h85;
        8'h6A: galois_lookup_148 = 8'hFA;
        8'h6B: galois_lookup_148 = 8'h6E;
        8'h6C: galois_lookup_148 = 8'h04;
        8'h6D: galois_lookup_148 = 8'h90;
        8'h6E: galois_lookup_148 = 8'hEF;
        8'h6F: galois_lookup_148 = 8'h7B;
        8'h70: galois_lookup_148 = 8'h6F;
        8'h71: galois_lookup_148 = 8'hFB;
        8'h72: galois_lookup_148 = 8'h84;
        8'h73: galois_lookup_148 = 8'h10;
        8'h74: galois_lookup_148 = 8'h7A;
        8'h75: galois_lookup_148 = 8'hEE;
        8'h76: galois_lookup_148 = 8'h91;
        8'h77: galois_lookup_148 = 8'h05;
        8'h78: galois_lookup_148 = 8'h45;
        8'h79: galois_lookup_148 = 8'hD1;
        8'h7A: galois_lookup_148 = 8'hAE;
        8'h7B: galois_lookup_148 = 8'h3A;
        8'h7C: galois_lookup_148 = 8'h50;
        8'h7D: galois_lookup_148 = 8'hC4;
        8'h7E: galois_lookup_148 = 8'hBB;
        8'h7F: galois_lookup_148 = 8'h2F;
        8'h80: galois_lookup_148 = 8'hE5;
        8'h81: galois_lookup_148 = 8'h71;
        8'h82: galois_lookup_148 = 8'h0E;
        8'h83: galois_lookup_148 = 8'h9A;
        8'h84: galois_lookup_148 = 8'hF0;
        8'h85: galois_lookup_148 = 8'h64;
        8'h86: galois_lookup_148 = 8'h1B;
        8'h87: galois_lookup_148 = 8'h8F;
        8'h88: galois_lookup_148 = 8'hCF;
        8'h89: galois_lookup_148 = 8'h5B;
        8'h8A: galois_lookup_148 = 8'h24;
        8'h8B: galois_lookup_148 = 8'hB0;
        8'h8C: galois_lookup_148 = 8'hDA;
        8'h8D: galois_lookup_148 = 8'h4E;
        8'h8E: galois_lookup_148 = 8'h31;
        8'h8F: galois_lookup_148 = 8'hA5;
        8'h90: galois_lookup_148 = 8'hB1;
        8'h91: galois_lookup_148 = 8'h25;
        8'h92: galois_lookup_148 = 8'h5A;
        8'h93: galois_lookup_148 = 8'hCE;
        8'h94: galois_lookup_148 = 8'hA4;
        8'h95: galois_lookup_148 = 8'h30;
        8'h96: galois_lookup_148 = 8'h4F;
        8'h97: galois_lookup_148 = 8'hDB;
        8'h98: galois_lookup_148 = 8'h9B;
        8'h99: galois_lookup_148 = 8'h0F;
        8'h9A: galois_lookup_148 = 8'h70;
        8'h9B: galois_lookup_148 = 8'hE4;
        8'h9C: galois_lookup_148 = 8'h8E;
        8'h9D: galois_lookup_148 = 8'h1A;
        8'h9E: galois_lookup_148 = 8'h65;
        8'h9F: galois_lookup_148 = 8'hF1;
        8'hA0: galois_lookup_148 = 8'h4D;
        8'hA1: galois_lookup_148 = 8'hD9;
        8'hA2: galois_lookup_148 = 8'hA6;
        8'hA3: galois_lookup_148 = 8'h32;
        8'hA4: galois_lookup_148 = 8'h58;
        8'hA5: galois_lookup_148 = 8'hCC;
        8'hA6: galois_lookup_148 = 8'hB3;
        8'hA7: galois_lookup_148 = 8'h27;
        8'hA8: galois_lookup_148 = 8'h67;
        8'hA9: galois_lookup_148 = 8'hF3;
        8'hAA: galois_lookup_148 = 8'h8C;
        8'hAB: galois_lookup_148 = 8'h18;
        8'hAC: galois_lookup_148 = 8'h72;
        8'hAD: galois_lookup_148 = 8'hE6;
        8'hAE: galois_lookup_148 = 8'h99;
        8'hAF: galois_lookup_148 = 8'h0D;
        8'hB0: galois_lookup_148 = 8'h19;
        8'hB1: galois_lookup_148 = 8'h8D;
        8'hB2: galois_lookup_148 = 8'hF2;
        8'hB3: galois_lookup_148 = 8'h66;
        8'hB4: galois_lookup_148 = 8'h0C;
        8'hB5: galois_lookup_148 = 8'h98;
        8'hB6: galois_lookup_148 = 8'hE7;
        8'hB7: galois_lookup_148 = 8'h73;
        8'hB8: galois_lookup_148 = 8'h33;
        8'hB9: galois_lookup_148 = 8'hA7;
        8'hBA: galois_lookup_148 = 8'hD8;
        8'hBB: galois_lookup_148 = 8'h4C;
        8'hBC: galois_lookup_148 = 8'h26;
        8'hBD: galois_lookup_148 = 8'hB2;
        8'hBE: galois_lookup_148 = 8'hCD;
        8'hBF: galois_lookup_148 = 8'h59;
        8'hC0: galois_lookup_148 = 8'h76;
        8'hC1: galois_lookup_148 = 8'hE2;
        8'hC2: galois_lookup_148 = 8'h9D;
        8'hC3: galois_lookup_148 = 8'h09;
        8'hC4: galois_lookup_148 = 8'h63;
        8'hC5: galois_lookup_148 = 8'hF7;
        8'hC6: galois_lookup_148 = 8'h88;
        8'hC7: galois_lookup_148 = 8'h1C;
        8'hC8: galois_lookup_148 = 8'h5C;
        8'hC9: galois_lookup_148 = 8'hC8;
        8'hCA: galois_lookup_148 = 8'hB7;
        8'hCB: galois_lookup_148 = 8'h23;
        8'hCC: galois_lookup_148 = 8'h49;
        8'hCD: galois_lookup_148 = 8'hDD;
        8'hCE: galois_lookup_148 = 8'hA2;
        8'hCF: galois_lookup_148 = 8'h36;
        8'hD0: galois_lookup_148 = 8'h22;
        8'hD1: galois_lookup_148 = 8'hB6;
        8'hD2: galois_lookup_148 = 8'hC9;
        8'hD3: galois_lookup_148 = 8'h5D;
        8'hD4: galois_lookup_148 = 8'h37;
        8'hD5: galois_lookup_148 = 8'hA3;
        8'hD6: galois_lookup_148 = 8'hDC;
        8'hD7: galois_lookup_148 = 8'h48;
        8'hD8: galois_lookup_148 = 8'h08;
        8'hD9: galois_lookup_148 = 8'h9C;
        8'hDA: galois_lookup_148 = 8'hE3;
        8'hDB: galois_lookup_148 = 8'h77;
        8'hDC: galois_lookup_148 = 8'h1D;
        8'hDD: galois_lookup_148 = 8'h89;
        8'hDE: galois_lookup_148 = 8'hF6;
        8'hDF: galois_lookup_148 = 8'h62;
        8'hE0: galois_lookup_148 = 8'hDE;
        8'hE1: galois_lookup_148 = 8'h4A;
        8'hE2: galois_lookup_148 = 8'h35;
        8'hE3: galois_lookup_148 = 8'hA1;
        8'hE4: galois_lookup_148 = 8'hCB;
        8'hE5: galois_lookup_148 = 8'h5F;
        8'hE6: galois_lookup_148 = 8'h20;
        8'hE7: galois_lookup_148 = 8'hB4;
        8'hE8: galois_lookup_148 = 8'hF4;
        8'hE9: galois_lookup_148 = 8'h60;
        8'hEA: galois_lookup_148 = 8'h1F;
        8'hEB: galois_lookup_148 = 8'h8B;
        8'hEC: galois_lookup_148 = 8'hE1;
        8'hED: galois_lookup_148 = 8'h75;
        8'hEE: galois_lookup_148 = 8'h0A;
        8'hEF: galois_lookup_148 = 8'h9E;
        8'hF0: galois_lookup_148 = 8'h8A;
        8'hF1: galois_lookup_148 = 8'h1E;
        8'hF2: galois_lookup_148 = 8'h61;
        8'hF3: galois_lookup_148 = 8'hF5;
        8'hF4: galois_lookup_148 = 8'h9F;
        8'hF5: galois_lookup_148 = 8'h0B;
        8'hF6: galois_lookup_148 = 8'h74;
        8'hF7: galois_lookup_148 = 8'hE0;
        8'hF8: galois_lookup_148 = 8'hA0;
        8'hF9: galois_lookup_148 = 8'h34;
        8'hFA: galois_lookup_148 = 8'h4B;
        8'hFB: galois_lookup_148 = 8'hDF;
        8'hFC: galois_lookup_148 = 8'hB5;
        8'hFD: galois_lookup_148 = 8'h21;
        8'hFE: galois_lookup_148 = 8'h5E;
        8'hFF: galois_lookup_148 = 8'hCA;
    endcase end
endfunction

// -----------------------------------------------------------------------------
function automatic [7:0] galois_lookup_192;
/*

*/
    input   [7:0]   byte;

    begin case (byte)
        8'h00: galois_lookup_192 = 8'h00;
        8'h01: galois_lookup_192 = 8'hC0;
        8'h02: galois_lookup_192 = 8'h43;
        8'h03: galois_lookup_192 = 8'h83;
        8'h04: galois_lookup_192 = 8'h86;
        8'h05: galois_lookup_192 = 8'h46;
        8'h06: galois_lookup_192 = 8'hC5;
        8'h07: galois_lookup_192 = 8'h05;
        8'h08: galois_lookup_192 = 8'hCF;
        8'h09: galois_lookup_192 = 8'h0F;
        8'h0A: galois_lookup_192 = 8'h8C;
        8'h0B: galois_lookup_192 = 8'h4C;
        8'h0C: galois_lookup_192 = 8'h49;
        8'h0D: galois_lookup_192 = 8'h89;
        8'h0E: galois_lookup_192 = 8'h0A;
        8'h0F: galois_lookup_192 = 8'hCA;
        8'h10: galois_lookup_192 = 8'h5D;
        8'h11: galois_lookup_192 = 8'h9D;
        8'h12: galois_lookup_192 = 8'h1E;
        8'h13: galois_lookup_192 = 8'hDE;
        8'h14: galois_lookup_192 = 8'hDB;
        8'h15: galois_lookup_192 = 8'h1B;
        8'h16: galois_lookup_192 = 8'h98;
        8'h17: galois_lookup_192 = 8'h58;
        8'h18: galois_lookup_192 = 8'h92;
        8'h19: galois_lookup_192 = 8'h52;
        8'h1A: galois_lookup_192 = 8'hD1;
        8'h1B: galois_lookup_192 = 8'h11;
        8'h1C: galois_lookup_192 = 8'h14;
        8'h1D: galois_lookup_192 = 8'hD4;
        8'h1E: galois_lookup_192 = 8'h57;
        8'h1F: galois_lookup_192 = 8'h97;
        8'h20: galois_lookup_192 = 8'hBA;
        8'h21: galois_lookup_192 = 8'h7A;
        8'h22: galois_lookup_192 = 8'hF9;
        8'h23: galois_lookup_192 = 8'h39;
        8'h24: galois_lookup_192 = 8'h3C;
        8'h25: galois_lookup_192 = 8'hFC;
        8'h26: galois_lookup_192 = 8'h7F;
        8'h27: galois_lookup_192 = 8'hBF;
        8'h28: galois_lookup_192 = 8'h75;
        8'h29: galois_lookup_192 = 8'hB5;
        8'h2A: galois_lookup_192 = 8'h36;
        8'h2B: galois_lookup_192 = 8'hF6;
        8'h2C: galois_lookup_192 = 8'hF3;
        8'h2D: galois_lookup_192 = 8'h33;
        8'h2E: galois_lookup_192 = 8'hB0;
        8'h2F: galois_lookup_192 = 8'h70;
        8'h30: galois_lookup_192 = 8'hE7;
        8'h31: galois_lookup_192 = 8'h27;
        8'h32: galois_lookup_192 = 8'hA4;
        8'h33: galois_lookup_192 = 8'h64;
        8'h34: galois_lookup_192 = 8'h61;
        8'h35: galois_lookup_192 = 8'hA1;
        8'h36: galois_lookup_192 = 8'h22;
        8'h37: galois_lookup_192 = 8'hE2;
        8'h38: galois_lookup_192 = 8'h28;
        8'h39: galois_lookup_192 = 8'hE8;
        8'h3A: galois_lookup_192 = 8'h6B;
        8'h3B: galois_lookup_192 = 8'hAB;
        8'h3C: galois_lookup_192 = 8'hAE;
        8'h3D: galois_lookup_192 = 8'h6E;
        8'h3E: galois_lookup_192 = 8'hED;
        8'h3F: galois_lookup_192 = 8'h2D;
        8'h40: galois_lookup_192 = 8'hB7;
        8'h41: galois_lookup_192 = 8'h77;
        8'h42: galois_lookup_192 = 8'hF4;
        8'h43: galois_lookup_192 = 8'h34;
        8'h44: galois_lookup_192 = 8'h31;
        8'h45: galois_lookup_192 = 8'hF1;
        8'h46: galois_lookup_192 = 8'h72;
        8'h47: galois_lookup_192 = 8'hB2;
        8'h48: galois_lookup_192 = 8'h78;
        8'h49: galois_lookup_192 = 8'hB8;
        8'h4A: galois_lookup_192 = 8'h3B;
        8'h4B: galois_lookup_192 = 8'hFB;
        8'h4C: galois_lookup_192 = 8'hFE;
        8'h4D: galois_lookup_192 = 8'h3E;
        8'h4E: galois_lookup_192 = 8'hBD;
        8'h4F: galois_lookup_192 = 8'h7D;
        8'h50: galois_lookup_192 = 8'hEA;
        8'h51: galois_lookup_192 = 8'h2A;
        8'h52: galois_lookup_192 = 8'hA9;
        8'h53: galois_lookup_192 = 8'h69;
        8'h54: galois_lookup_192 = 8'h6C;
        8'h55: galois_lookup_192 = 8'hAC;
        8'h56: galois_lookup_192 = 8'h2F;
        8'h57: galois_lookup_192 = 8'hEF;
        8'h58: galois_lookup_192 = 8'h25;
        8'h59: galois_lookup_192 = 8'hE5;
        8'h5A: galois_lookup_192 = 8'h66;
        8'h5B: galois_lookup_192 = 8'hA6;
        8'h5C: galois_lookup_192 = 8'hA3;
        8'h5D: galois_lookup_192 = 8'h63;
        8'h5E: galois_lookup_192 = 8'hE0;
        8'h5F: galois_lookup_192 = 8'h20;
        8'h60: galois_lookup_192 = 8'h0D;
        8'h61: galois_lookup_192 = 8'hCD;
        8'h62: galois_lookup_192 = 8'h4E;
        8'h63: galois_lookup_192 = 8'h8E;
        8'h64: galois_lookup_192 = 8'h8B;
        8'h65: galois_lookup_192 = 8'h4B;
        8'h66: galois_lookup_192 = 8'hC8;
        8'h67: galois_lookup_192 = 8'h08;
        8'h68: galois_lookup_192 = 8'hC2;
        8'h69: galois_lookup_192 = 8'h02;
        8'h6A: galois_lookup_192 = 8'h81;
        8'h6B: galois_lookup_192 = 8'h41;
        8'h6C: galois_lookup_192 = 8'h44;
        8'h6D: galois_lookup_192 = 8'h84;
        8'h6E: galois_lookup_192 = 8'h07;
        8'h6F: galois_lookup_192 = 8'hC7;
        8'h70: galois_lookup_192 = 8'h50;
        8'h71: galois_lookup_192 = 8'h90;
        8'h72: galois_lookup_192 = 8'h13;
        8'h73: galois_lookup_192 = 8'hD3;
        8'h74: galois_lookup_192 = 8'hD6;
        8'h75: galois_lookup_192 = 8'h16;
        8'h76: galois_lookup_192 = 8'h95;
        8'h77: galois_lookup_192 = 8'h55;
        8'h78: galois_lookup_192 = 8'h9F;
        8'h79: galois_lookup_192 = 8'h5F;
        8'h7A: galois_lookup_192 = 8'hDC;
        8'h7B: galois_lookup_192 = 8'h1C;
        8'h7C: galois_lookup_192 = 8'h19;
        8'h7D: galois_lookup_192 = 8'hD9;
        8'h7E: galois_lookup_192 = 8'h5A;
        8'h7F: galois_lookup_192 = 8'h9A;
        8'h80: galois_lookup_192 = 8'hAD;
        8'h81: galois_lookup_192 = 8'h6D;
        8'h82: galois_lookup_192 = 8'hEE;
        8'h83: galois_lookup_192 = 8'h2E;
        8'h84: galois_lookup_192 = 8'h2B;
        8'h85: galois_lookup_192 = 8'hEB;
        8'h86: galois_lookup_192 = 8'h68;
        8'h87: galois_lookup_192 = 8'hA8;
        8'h88: galois_lookup_192 = 8'h62;
        8'h89: galois_lookup_192 = 8'hA2;
        8'h8A: galois_lookup_192 = 8'h21;
        8'h8B: galois_lookup_192 = 8'hE1;
        8'h8C: galois_lookup_192 = 8'hE4;
        8'h8D: galois_lookup_192 = 8'h24;
        8'h8E: galois_lookup_192 = 8'hA7;
        8'h8F: galois_lookup_192 = 8'h67;
        8'h90: galois_lookup_192 = 8'hF0;
        8'h91: galois_lookup_192 = 8'h30;
        8'h92: galois_lookup_192 = 8'hB3;
        8'h93: galois_lookup_192 = 8'h73;
        8'h94: galois_lookup_192 = 8'h76;
        8'h95: galois_lookup_192 = 8'hB6;
        8'h96: galois_lookup_192 = 8'h35;
        8'h97: galois_lookup_192 = 8'hF5;
        8'h98: galois_lookup_192 = 8'h3F;
        8'h99: galois_lookup_192 = 8'hFF;
        8'h9A: galois_lookup_192 = 8'h7C;
        8'h9B: galois_lookup_192 = 8'hBC;
        8'h9C: galois_lookup_192 = 8'hB9;
        8'h9D: galois_lookup_192 = 8'h79;
        8'h9E: galois_lookup_192 = 8'hFA;
        8'h9F: galois_lookup_192 = 8'h3A;
        8'hA0: galois_lookup_192 = 8'h17;
        8'hA1: galois_lookup_192 = 8'hD7;
        8'hA2: galois_lookup_192 = 8'h54;
        8'hA3: galois_lookup_192 = 8'h94;
        8'hA4: galois_lookup_192 = 8'h91;
        8'hA5: galois_lookup_192 = 8'h51;
        8'hA6: galois_lookup_192 = 8'hD2;
        8'hA7: galois_lookup_192 = 8'h12;
        8'hA8: galois_lookup_192 = 8'hD8;
        8'hA9: galois_lookup_192 = 8'h18;
        8'hAA: galois_lookup_192 = 8'h9B;
        8'hAB: galois_lookup_192 = 8'h5B;
        8'hAC: galois_lookup_192 = 8'h5E;
        8'hAD: galois_lookup_192 = 8'h9E;
        8'hAE: galois_lookup_192 = 8'h1D;
        8'hAF: galois_lookup_192 = 8'hDD;
        8'hB0: galois_lookup_192 = 8'h4A;
        8'hB1: galois_lookup_192 = 8'h8A;
        8'hB2: galois_lookup_192 = 8'h09;
        8'hB3: galois_lookup_192 = 8'hC9;
        8'hB4: galois_lookup_192 = 8'hCC;
        8'hB5: galois_lookup_192 = 8'h0C;
        8'hB6: galois_lookup_192 = 8'h8F;
        8'hB7: galois_lookup_192 = 8'h4F;
        8'hB8: galois_lookup_192 = 8'h85;
        8'hB9: galois_lookup_192 = 8'h45;
        8'hBA: galois_lookup_192 = 8'hC6;
        8'hBB: galois_lookup_192 = 8'h06;
        8'hBC: galois_lookup_192 = 8'h03;
        8'hBD: galois_lookup_192 = 8'hC3;
        8'hBE: galois_lookup_192 = 8'h40;
        8'hBF: galois_lookup_192 = 8'h80;
        8'hC0: galois_lookup_192 = 8'h1A;
        8'hC1: galois_lookup_192 = 8'hDA;
        8'hC2: galois_lookup_192 = 8'h59;
        8'hC3: galois_lookup_192 = 8'h99;
        8'hC4: galois_lookup_192 = 8'h9C;
        8'hC5: galois_lookup_192 = 8'h5C;
        8'hC6: galois_lookup_192 = 8'hDF;
        8'hC7: galois_lookup_192 = 8'h1F;
        8'hC8: galois_lookup_192 = 8'hD5;
        8'hC9: galois_lookup_192 = 8'h15;
        8'hCA: galois_lookup_192 = 8'h96;
        8'hCB: galois_lookup_192 = 8'h56;
        8'hCC: galois_lookup_192 = 8'h53;
        8'hCD: galois_lookup_192 = 8'h93;
        8'hCE: galois_lookup_192 = 8'h10;
        8'hCF: galois_lookup_192 = 8'hD0;
        8'hD0: galois_lookup_192 = 8'h47;
        8'hD1: galois_lookup_192 = 8'h87;
        8'hD2: galois_lookup_192 = 8'h04;
        8'hD3: galois_lookup_192 = 8'hC4;
        8'hD4: galois_lookup_192 = 8'hC1;
        8'hD5: galois_lookup_192 = 8'h01;
        8'hD6: galois_lookup_192 = 8'h82;
        8'hD7: galois_lookup_192 = 8'h42;
        8'hD8: galois_lookup_192 = 8'h88;
        8'hD9: galois_lookup_192 = 8'h48;
        8'hDA: galois_lookup_192 = 8'hCB;
        8'hDB: galois_lookup_192 = 8'h0B;
        8'hDC: galois_lookup_192 = 8'h0E;
        8'hDD: galois_lookup_192 = 8'hCE;
        8'hDE: galois_lookup_192 = 8'h4D;
        8'hDF: galois_lookup_192 = 8'h8D;
        8'hE0: galois_lookup_192 = 8'hA0;
        8'hE1: galois_lookup_192 = 8'h60;
        8'hE2: galois_lookup_192 = 8'hE3;
        8'hE3: galois_lookup_192 = 8'h23;
        8'hE4: galois_lookup_192 = 8'h26;
        8'hE5: galois_lookup_192 = 8'hE6;
        8'hE6: galois_lookup_192 = 8'h65;
        8'hE7: galois_lookup_192 = 8'hA5;
        8'hE8: galois_lookup_192 = 8'h6F;
        8'hE9: galois_lookup_192 = 8'hAF;
        8'hEA: galois_lookup_192 = 8'h2C;
        8'hEB: galois_lookup_192 = 8'hEC;
        8'hEC: galois_lookup_192 = 8'hE9;
        8'hED: galois_lookup_192 = 8'h29;
        8'hEE: galois_lookup_192 = 8'hAA;
        8'hEF: galois_lookup_192 = 8'h6A;
        8'hF0: galois_lookup_192 = 8'hFD;
        8'hF1: galois_lookup_192 = 8'h3D;
        8'hF2: galois_lookup_192 = 8'hBE;
        8'hF3: galois_lookup_192 = 8'h7E;
        8'hF4: galois_lookup_192 = 8'h7B;
        8'hF5: galois_lookup_192 = 8'hBB;
        8'hF6: galois_lookup_192 = 8'h38;
        8'hF7: galois_lookup_192 = 8'hF8;
        8'hF8: galois_lookup_192 = 8'h32;
        8'hF9: galois_lookup_192 = 8'hF2;
        8'hFA: galois_lookup_192 = 8'h71;
        8'hFB: galois_lookup_192 = 8'hB1;
        8'hFC: galois_lookup_192 = 8'hB4;
        8'hFD: galois_lookup_192 = 8'h74;
        8'hFE: galois_lookup_192 = 8'hF7;
        8'hFF: galois_lookup_192 = 8'h37;
    endcase end
endfunction

// -----------------------------------------------------------------------------
function automatic [7:0] galois_lookup_194;
/*

*/
    input   [7:0]   byte;

    begin case (byte)
        8'h00: galois_lookup_194 = 8'h00;
        8'h01: galois_lookup_194 = 8'hC2;
        8'h02: galois_lookup_194 = 8'h47;
        8'h03: galois_lookup_194 = 8'h85;
        8'h04: galois_lookup_194 = 8'h8E;
        8'h05: galois_lookup_194 = 8'h4C;
        8'h06: galois_lookup_194 = 8'hC9;
        8'h07: galois_lookup_194 = 8'h0B;
        8'h08: galois_lookup_194 = 8'hDF;
        8'h09: galois_lookup_194 = 8'h1D;
        8'h0A: galois_lookup_194 = 8'h98;
        8'h0B: galois_lookup_194 = 8'h5A;
        8'h0C: galois_lookup_194 = 8'h51;
        8'h0D: galois_lookup_194 = 8'h93;
        8'h0E: galois_lookup_194 = 8'h16;
        8'h0F: galois_lookup_194 = 8'hD4;
        8'h10: galois_lookup_194 = 8'h7D;
        8'h11: galois_lookup_194 = 8'hBF;
        8'h12: galois_lookup_194 = 8'h3A;
        8'h13: galois_lookup_194 = 8'hF8;
        8'h14: galois_lookup_194 = 8'hF3;
        8'h15: galois_lookup_194 = 8'h31;
        8'h16: galois_lookup_194 = 8'hB4;
        8'h17: galois_lookup_194 = 8'h76;
        8'h18: galois_lookup_194 = 8'hA2;
        8'h19: galois_lookup_194 = 8'h60;
        8'h1A: galois_lookup_194 = 8'hE5;
        8'h1B: galois_lookup_194 = 8'h27;
        8'h1C: galois_lookup_194 = 8'h2C;
        8'h1D: galois_lookup_194 = 8'hEE;
        8'h1E: galois_lookup_194 = 8'h6B;
        8'h1F: galois_lookup_194 = 8'hA9;
        8'h20: galois_lookup_194 = 8'hFA;
        8'h21: galois_lookup_194 = 8'h38;
        8'h22: galois_lookup_194 = 8'hBD;
        8'h23: galois_lookup_194 = 8'h7F;
        8'h24: galois_lookup_194 = 8'h74;
        8'h25: galois_lookup_194 = 8'hB6;
        8'h26: galois_lookup_194 = 8'h33;
        8'h27: galois_lookup_194 = 8'hF1;
        8'h28: galois_lookup_194 = 8'h25;
        8'h29: galois_lookup_194 = 8'hE7;
        8'h2A: galois_lookup_194 = 8'h62;
        8'h2B: galois_lookup_194 = 8'hA0;
        8'h2C: galois_lookup_194 = 8'hAB;
        8'h2D: galois_lookup_194 = 8'h69;
        8'h2E: galois_lookup_194 = 8'hEC;
        8'h2F: galois_lookup_194 = 8'h2E;
        8'h30: galois_lookup_194 = 8'h87;
        8'h31: galois_lookup_194 = 8'h45;
        8'h32: galois_lookup_194 = 8'hC0;
        8'h33: galois_lookup_194 = 8'h02;
        8'h34: galois_lookup_194 = 8'h09;
        8'h35: galois_lookup_194 = 8'hCB;
        8'h36: galois_lookup_194 = 8'h4E;
        8'h37: galois_lookup_194 = 8'h8C;
        8'h38: galois_lookup_194 = 8'h58;
        8'h39: galois_lookup_194 = 8'h9A;
        8'h3A: galois_lookup_194 = 8'h1F;
        8'h3B: galois_lookup_194 = 8'hDD;
        8'h3C: galois_lookup_194 = 8'hD6;
        8'h3D: galois_lookup_194 = 8'h14;
        8'h3E: galois_lookup_194 = 8'h91;
        8'h3F: galois_lookup_194 = 8'h53;
        8'h40: galois_lookup_194 = 8'h37;
        8'h41: galois_lookup_194 = 8'hF5;
        8'h42: galois_lookup_194 = 8'h70;
        8'h43: galois_lookup_194 = 8'hB2;
        8'h44: galois_lookup_194 = 8'hB9;
        8'h45: galois_lookup_194 = 8'h7B;
        8'h46: galois_lookup_194 = 8'hFE;
        8'h47: galois_lookup_194 = 8'h3C;
        8'h48: galois_lookup_194 = 8'hE8;
        8'h49: galois_lookup_194 = 8'h2A;
        8'h4A: galois_lookup_194 = 8'hAF;
        8'h4B: galois_lookup_194 = 8'h6D;
        8'h4C: galois_lookup_194 = 8'h66;
        8'h4D: galois_lookup_194 = 8'hA4;
        8'h4E: galois_lookup_194 = 8'h21;
        8'h4F: galois_lookup_194 = 8'hE3;
        8'h50: galois_lookup_194 = 8'h4A;
        8'h51: galois_lookup_194 = 8'h88;
        8'h52: galois_lookup_194 = 8'h0D;
        8'h53: galois_lookup_194 = 8'hCF;
        8'h54: galois_lookup_194 = 8'hC4;
        8'h55: galois_lookup_194 = 8'h06;
        8'h56: galois_lookup_194 = 8'h83;
        8'h57: galois_lookup_194 = 8'h41;
        8'h58: galois_lookup_194 = 8'h95;
        8'h59: galois_lookup_194 = 8'h57;
        8'h5A: galois_lookup_194 = 8'hD2;
        8'h5B: galois_lookup_194 = 8'h10;
        8'h5C: galois_lookup_194 = 8'h1B;
        8'h5D: galois_lookup_194 = 8'hD9;
        8'h5E: galois_lookup_194 = 8'h5C;
        8'h5F: galois_lookup_194 = 8'h9E;
        8'h60: galois_lookup_194 = 8'hCD;
        8'h61: galois_lookup_194 = 8'h0F;
        8'h62: galois_lookup_194 = 8'h8A;
        8'h63: galois_lookup_194 = 8'h48;
        8'h64: galois_lookup_194 = 8'h43;
        8'h65: galois_lookup_194 = 8'h81;
        8'h66: galois_lookup_194 = 8'h04;
        8'h67: galois_lookup_194 = 8'hC6;
        8'h68: galois_lookup_194 = 8'h12;
        8'h69: galois_lookup_194 = 8'hD0;
        8'h6A: galois_lookup_194 = 8'h55;
        8'h6B: galois_lookup_194 = 8'h97;
        8'h6C: galois_lookup_194 = 8'h9C;
        8'h6D: galois_lookup_194 = 8'h5E;
        8'h6E: galois_lookup_194 = 8'hDB;
        8'h6F: galois_lookup_194 = 8'h19;
        8'h70: galois_lookup_194 = 8'hB0;
        8'h71: galois_lookup_194 = 8'h72;
        8'h72: galois_lookup_194 = 8'hF7;
        8'h73: galois_lookup_194 = 8'h35;
        8'h74: galois_lookup_194 = 8'h3E;
        8'h75: galois_lookup_194 = 8'hFC;
        8'h76: galois_lookup_194 = 8'h79;
        8'h77: galois_lookup_194 = 8'hBB;
        8'h78: galois_lookup_194 = 8'h6F;
        8'h79: galois_lookup_194 = 8'hAD;
        8'h7A: galois_lookup_194 = 8'h28;
        8'h7B: galois_lookup_194 = 8'hEA;
        8'h7C: galois_lookup_194 = 8'hE1;
        8'h7D: galois_lookup_194 = 8'h23;
        8'h7E: galois_lookup_194 = 8'hA6;
        8'h7F: galois_lookup_194 = 8'h64;
        8'h80: galois_lookup_194 = 8'h6E;
        8'h81: galois_lookup_194 = 8'hAC;
        8'h82: galois_lookup_194 = 8'h29;
        8'h83: galois_lookup_194 = 8'hEB;
        8'h84: galois_lookup_194 = 8'hE0;
        8'h85: galois_lookup_194 = 8'h22;
        8'h86: galois_lookup_194 = 8'hA7;
        8'h87: galois_lookup_194 = 8'h65;
        8'h88: galois_lookup_194 = 8'hB1;
        8'h89: galois_lookup_194 = 8'h73;
        8'h8A: galois_lookup_194 = 8'hF6;
        8'h8B: galois_lookup_194 = 8'h34;
        8'h8C: galois_lookup_194 = 8'h3F;
        8'h8D: galois_lookup_194 = 8'hFD;
        8'h8E: galois_lookup_194 = 8'h78;
        8'h8F: galois_lookup_194 = 8'hBA;
        8'h90: galois_lookup_194 = 8'h13;
        8'h91: galois_lookup_194 = 8'hD1;
        8'h92: galois_lookup_194 = 8'h54;
        8'h93: galois_lookup_194 = 8'h96;
        8'h94: galois_lookup_194 = 8'h9D;
        8'h95: galois_lookup_194 = 8'h5F;
        8'h96: galois_lookup_194 = 8'hDA;
        8'h97: galois_lookup_194 = 8'h18;
        8'h98: galois_lookup_194 = 8'hCC;
        8'h99: galois_lookup_194 = 8'h0E;
        8'h9A: galois_lookup_194 = 8'h8B;
        8'h9B: galois_lookup_194 = 8'h49;
        8'h9C: galois_lookup_194 = 8'h42;
        8'h9D: galois_lookup_194 = 8'h80;
        8'h9E: galois_lookup_194 = 8'h05;
        8'h9F: galois_lookup_194 = 8'hC7;
        8'hA0: galois_lookup_194 = 8'h94;
        8'hA1: galois_lookup_194 = 8'h56;
        8'hA2: galois_lookup_194 = 8'hD3;
        8'hA3: galois_lookup_194 = 8'h11;
        8'hA4: galois_lookup_194 = 8'h1A;
        8'hA5: galois_lookup_194 = 8'hD8;
        8'hA6: galois_lookup_194 = 8'h5D;
        8'hA7: galois_lookup_194 = 8'h9F;
        8'hA8: galois_lookup_194 = 8'h4B;
        8'hA9: galois_lookup_194 = 8'h89;
        8'hAA: galois_lookup_194 = 8'h0C;
        8'hAB: galois_lookup_194 = 8'hCE;
        8'hAC: galois_lookup_194 = 8'hC5;
        8'hAD: galois_lookup_194 = 8'h07;
        8'hAE: galois_lookup_194 = 8'h82;
        8'hAF: galois_lookup_194 = 8'h40;
        8'hB0: galois_lookup_194 = 8'hE9;
        8'hB1: galois_lookup_194 = 8'h2B;
        8'hB2: galois_lookup_194 = 8'hAE;
        8'hB3: galois_lookup_194 = 8'h6C;
        8'hB4: galois_lookup_194 = 8'h67;
        8'hB5: galois_lookup_194 = 8'hA5;
        8'hB6: galois_lookup_194 = 8'h20;
        8'hB7: galois_lookup_194 = 8'hE2;
        8'hB8: galois_lookup_194 = 8'h36;
        8'hB9: galois_lookup_194 = 8'hF4;
        8'hBA: galois_lookup_194 = 8'h71;
        8'hBB: galois_lookup_194 = 8'hB3;
        8'hBC: galois_lookup_194 = 8'hB8;
        8'hBD: galois_lookup_194 = 8'h7A;
        8'hBE: galois_lookup_194 = 8'hFF;
        8'hBF: galois_lookup_194 = 8'h3D;
        8'hC0: galois_lookup_194 = 8'h59;
        8'hC1: galois_lookup_194 = 8'h9B;
        8'hC2: galois_lookup_194 = 8'h1E;
        8'hC3: galois_lookup_194 = 8'hDC;
        8'hC4: galois_lookup_194 = 8'hD7;
        8'hC5: galois_lookup_194 = 8'h15;
        8'hC6: galois_lookup_194 = 8'h90;
        8'hC7: galois_lookup_194 = 8'h52;
        8'hC8: galois_lookup_194 = 8'h86;
        8'hC9: galois_lookup_194 = 8'h44;
        8'hCA: galois_lookup_194 = 8'hC1;
        8'hCB: galois_lookup_194 = 8'h03;
        8'hCC: galois_lookup_194 = 8'h08;
        8'hCD: galois_lookup_194 = 8'hCA;
        8'hCE: galois_lookup_194 = 8'h4F;
        8'hCF: galois_lookup_194 = 8'h8D;
        8'hD0: galois_lookup_194 = 8'h24;
        8'hD1: galois_lookup_194 = 8'hE6;
        8'hD2: galois_lookup_194 = 8'h63;
        8'hD3: galois_lookup_194 = 8'hA1;
        8'hD4: galois_lookup_194 = 8'hAA;
        8'hD5: galois_lookup_194 = 8'h68;
        8'hD6: galois_lookup_194 = 8'hED;
        8'hD7: galois_lookup_194 = 8'h2F;
        8'hD8: galois_lookup_194 = 8'hFB;
        8'hD9: galois_lookup_194 = 8'h39;
        8'hDA: galois_lookup_194 = 8'hBC;
        8'hDB: galois_lookup_194 = 8'h7E;
        8'hDC: galois_lookup_194 = 8'h75;
        8'hDD: galois_lookup_194 = 8'hB7;
        8'hDE: galois_lookup_194 = 8'h32;
        8'hDF: galois_lookup_194 = 8'hF0;
        8'hE0: galois_lookup_194 = 8'hA3;
        8'hE1: galois_lookup_194 = 8'h61;
        8'hE2: galois_lookup_194 = 8'hE4;
        8'hE3: galois_lookup_194 = 8'h26;
        8'hE4: galois_lookup_194 = 8'h2D;
        8'hE5: galois_lookup_194 = 8'hEF;
        8'hE6: galois_lookup_194 = 8'h6A;
        8'hE7: galois_lookup_194 = 8'hA8;
        8'hE8: galois_lookup_194 = 8'h7C;
        8'hE9: galois_lookup_194 = 8'hBE;
        8'hEA: galois_lookup_194 = 8'h3B;
        8'hEB: galois_lookup_194 = 8'hF9;
        8'hEC: galois_lookup_194 = 8'hF2;
        8'hED: galois_lookup_194 = 8'h30;
        8'hEE: galois_lookup_194 = 8'hB5;
        8'hEF: galois_lookup_194 = 8'h77;
        8'hF0: galois_lookup_194 = 8'hDE;
        8'hF1: galois_lookup_194 = 8'h1C;
        8'hF2: galois_lookup_194 = 8'h99;
        8'hF3: galois_lookup_194 = 8'h5B;
        8'hF4: galois_lookup_194 = 8'h50;
        8'hF5: galois_lookup_194 = 8'h92;
        8'hF6: galois_lookup_194 = 8'h17;
        8'hF7: galois_lookup_194 = 8'hD5;
        8'hF8: galois_lookup_194 = 8'h01;
        8'hF9: galois_lookup_194 = 8'hC3;
        8'hFA: galois_lookup_194 = 8'h46;
        8'hFB: galois_lookup_194 = 8'h84;
        8'hFC: galois_lookup_194 = 8'h8F;
        8'hFD: galois_lookup_194 = 8'h4D;
        8'hFE: galois_lookup_194 = 8'hC8;
        8'hFF: galois_lookup_194 = 8'h0A;
    endcase end
endfunction

// -----------------------------------------------------------------------------
function automatic [7:0] galois_lookup_251;
/*

*/
    input   [7:0]   byte;

    begin case (byte)
        8'h00: galois_lookup_251 = 8'h00;
        8'h01: galois_lookup_251 = 8'hFB;
        8'h02: galois_lookup_251 = 8'h35;
        8'h03: galois_lookup_251 = 8'hCE;
        8'h04: galois_lookup_251 = 8'h6A;
        8'h05: galois_lookup_251 = 8'h91;
        8'h06: galois_lookup_251 = 8'h5F;
        8'h07: galois_lookup_251 = 8'hA4;
        8'h08: galois_lookup_251 = 8'hD4;
        8'h09: galois_lookup_251 = 8'h2F;
        8'h0A: galois_lookup_251 = 8'hE1;
        8'h0B: galois_lookup_251 = 8'h1A;
        8'h0C: galois_lookup_251 = 8'hBE;
        8'h0D: galois_lookup_251 = 8'h45;
        8'h0E: galois_lookup_251 = 8'h8B;
        8'h0F: galois_lookup_251 = 8'h70;
        8'h10: galois_lookup_251 = 8'h6B;
        8'h11: galois_lookup_251 = 8'h90;
        8'h12: galois_lookup_251 = 8'h5E;
        8'h13: galois_lookup_251 = 8'hA5;
        8'h14: galois_lookup_251 = 8'h01;
        8'h15: galois_lookup_251 = 8'hFA;
        8'h16: galois_lookup_251 = 8'h34;
        8'h17: galois_lookup_251 = 8'hCF;
        8'h18: galois_lookup_251 = 8'hBF;
        8'h19: galois_lookup_251 = 8'h44;
        8'h1A: galois_lookup_251 = 8'h8A;
        8'h1B: galois_lookup_251 = 8'h71;
        8'h1C: galois_lookup_251 = 8'hD5;
        8'h1D: galois_lookup_251 = 8'h2E;
        8'h1E: galois_lookup_251 = 8'hE0;
        8'h1F: galois_lookup_251 = 8'h1B;
        8'h20: galois_lookup_251 = 8'hD6;
        8'h21: galois_lookup_251 = 8'h2D;
        8'h22: galois_lookup_251 = 8'hE3;
        8'h23: galois_lookup_251 = 8'h18;
        8'h24: galois_lookup_251 = 8'hBC;
        8'h25: galois_lookup_251 = 8'h47;
        8'h26: galois_lookup_251 = 8'h89;
        8'h27: galois_lookup_251 = 8'h72;
        8'h28: galois_lookup_251 = 8'h02;
        8'h29: galois_lookup_251 = 8'hF9;
        8'h2A: galois_lookup_251 = 8'h37;
        8'h2B: galois_lookup_251 = 8'hCC;
        8'h2C: galois_lookup_251 = 8'h68;
        8'h2D: galois_lookup_251 = 8'h93;
        8'h2E: galois_lookup_251 = 8'h5D;
        8'h2F: galois_lookup_251 = 8'hA6;
        8'h30: galois_lookup_251 = 8'hBD;
        8'h31: galois_lookup_251 = 8'h46;
        8'h32: galois_lookup_251 = 8'h88;
        8'h33: galois_lookup_251 = 8'h73;
        8'h34: galois_lookup_251 = 8'hD7;
        8'h35: galois_lookup_251 = 8'h2C;
        8'h36: galois_lookup_251 = 8'hE2;
        8'h37: galois_lookup_251 = 8'h19;
        8'h38: galois_lookup_251 = 8'h69;
        8'h39: galois_lookup_251 = 8'h92;
        8'h3A: galois_lookup_251 = 8'h5C;
        8'h3B: galois_lookup_251 = 8'hA7;
        8'h3C: galois_lookup_251 = 8'h03;
        8'h3D: galois_lookup_251 = 8'hF8;
        8'h3E: galois_lookup_251 = 8'h36;
        8'h3F: galois_lookup_251 = 8'hCD;
        8'h40: galois_lookup_251 = 8'h6F;
        8'h41: galois_lookup_251 = 8'h94;
        8'h42: galois_lookup_251 = 8'h5A;
        8'h43: galois_lookup_251 = 8'hA1;
        8'h44: galois_lookup_251 = 8'h05;
        8'h45: galois_lookup_251 = 8'hFE;
        8'h46: galois_lookup_251 = 8'h30;
        8'h47: galois_lookup_251 = 8'hCB;
        8'h48: galois_lookup_251 = 8'hBB;
        8'h49: galois_lookup_251 = 8'h40;
        8'h4A: galois_lookup_251 = 8'h8E;
        8'h4B: galois_lookup_251 = 8'h75;
        8'h4C: galois_lookup_251 = 8'hD1;
        8'h4D: galois_lookup_251 = 8'h2A;
        8'h4E: galois_lookup_251 = 8'hE4;
        8'h4F: galois_lookup_251 = 8'h1F;
        8'h50: galois_lookup_251 = 8'h04;
        8'h51: galois_lookup_251 = 8'hFF;
        8'h52: galois_lookup_251 = 8'h31;
        8'h53: galois_lookup_251 = 8'hCA;
        8'h54: galois_lookup_251 = 8'h6E;
        8'h55: galois_lookup_251 = 8'h95;
        8'h56: galois_lookup_251 = 8'h5B;
        8'h57: galois_lookup_251 = 8'hA0;
        8'h58: galois_lookup_251 = 8'hD0;
        8'h59: galois_lookup_251 = 8'h2B;
        8'h5A: galois_lookup_251 = 8'hE5;
        8'h5B: galois_lookup_251 = 8'h1E;
        8'h5C: galois_lookup_251 = 8'hBA;
        8'h5D: galois_lookup_251 = 8'h41;
        8'h5E: galois_lookup_251 = 8'h8F;
        8'h5F: galois_lookup_251 = 8'h74;
        8'h60: galois_lookup_251 = 8'hB9;
        8'h61: galois_lookup_251 = 8'h42;
        8'h62: galois_lookup_251 = 8'h8C;
        8'h63: galois_lookup_251 = 8'h77;
        8'h64: galois_lookup_251 = 8'hD3;
        8'h65: galois_lookup_251 = 8'h28;
        8'h66: galois_lookup_251 = 8'hE6;
        8'h67: galois_lookup_251 = 8'h1D;
        8'h68: galois_lookup_251 = 8'h6D;
        8'h69: galois_lookup_251 = 8'h96;
        8'h6A: galois_lookup_251 = 8'h58;
        8'h6B: galois_lookup_251 = 8'hA3;
        8'h6C: galois_lookup_251 = 8'h07;
        8'h6D: galois_lookup_251 = 8'hFC;
        8'h6E: galois_lookup_251 = 8'h32;
        8'h6F: galois_lookup_251 = 8'hC9;
        8'h70: galois_lookup_251 = 8'hD2;
        8'h71: galois_lookup_251 = 8'h29;
        8'h72: galois_lookup_251 = 8'hE7;
        8'h73: galois_lookup_251 = 8'h1C;
        8'h74: galois_lookup_251 = 8'hB8;
        8'h75: galois_lookup_251 = 8'h43;
        8'h76: galois_lookup_251 = 8'h8D;
        8'h77: galois_lookup_251 = 8'h76;
        8'h78: galois_lookup_251 = 8'h06;
        8'h79: galois_lookup_251 = 8'hFD;
        8'h7A: galois_lookup_251 = 8'h33;
        8'h7B: galois_lookup_251 = 8'hC8;
        8'h7C: galois_lookup_251 = 8'h6C;
        8'h7D: galois_lookup_251 = 8'h97;
        8'h7E: galois_lookup_251 = 8'h59;
        8'h7F: galois_lookup_251 = 8'hA2;
        8'h80: galois_lookup_251 = 8'hDE;
        8'h81: galois_lookup_251 = 8'h25;
        8'h82: galois_lookup_251 = 8'hEB;
        8'h83: galois_lookup_251 = 8'h10;
        8'h84: galois_lookup_251 = 8'hB4;
        8'h85: galois_lookup_251 = 8'h4F;
        8'h86: galois_lookup_251 = 8'h81;
        8'h87: galois_lookup_251 = 8'h7A;
        8'h88: galois_lookup_251 = 8'h0A;
        8'h89: galois_lookup_251 = 8'hF1;
        8'h8A: galois_lookup_251 = 8'h3F;
        8'h8B: galois_lookup_251 = 8'hC4;
        8'h8C: galois_lookup_251 = 8'h60;
        8'h8D: galois_lookup_251 = 8'h9B;
        8'h8E: galois_lookup_251 = 8'h55;
        8'h8F: galois_lookup_251 = 8'hAE;
        8'h90: galois_lookup_251 = 8'hB5;
        8'h91: galois_lookup_251 = 8'h4E;
        8'h92: galois_lookup_251 = 8'h80;
        8'h93: galois_lookup_251 = 8'h7B;
        8'h94: galois_lookup_251 = 8'hDF;
        8'h95: galois_lookup_251 = 8'h24;
        8'h96: galois_lookup_251 = 8'hEA;
        8'h97: galois_lookup_251 = 8'h11;
        8'h98: galois_lookup_251 = 8'h61;
        8'h99: galois_lookup_251 = 8'h9A;
        8'h9A: galois_lookup_251 = 8'h54;
        8'h9B: galois_lookup_251 = 8'hAF;
        8'h9C: galois_lookup_251 = 8'h0B;
        8'h9D: galois_lookup_251 = 8'hF0;
        8'h9E: galois_lookup_251 = 8'h3E;
        8'h9F: galois_lookup_251 = 8'hC5;
        8'hA0: galois_lookup_251 = 8'h08;
        8'hA1: galois_lookup_251 = 8'hF3;
        8'hA2: galois_lookup_251 = 8'h3D;
        8'hA3: galois_lookup_251 = 8'hC6;
        8'hA4: galois_lookup_251 = 8'h62;
        8'hA5: galois_lookup_251 = 8'h99;
        8'hA6: galois_lookup_251 = 8'h57;
        8'hA7: galois_lookup_251 = 8'hAC;
        8'hA8: galois_lookup_251 = 8'hDC;
        8'hA9: galois_lookup_251 = 8'h27;
        8'hAA: galois_lookup_251 = 8'hE9;
        8'hAB: galois_lookup_251 = 8'h12;
        8'hAC: galois_lookup_251 = 8'hB6;
        8'hAD: galois_lookup_251 = 8'h4D;
        8'hAE: galois_lookup_251 = 8'h83;
        8'hAF: galois_lookup_251 = 8'h78;
        8'hB0: galois_lookup_251 = 8'h63;
        8'hB1: galois_lookup_251 = 8'h98;
        8'hB2: galois_lookup_251 = 8'h56;
        8'hB3: galois_lookup_251 = 8'hAD;
        8'hB4: galois_lookup_251 = 8'h09;
        8'hB5: galois_lookup_251 = 8'hF2;
        8'hB6: galois_lookup_251 = 8'h3C;
        8'hB7: galois_lookup_251 = 8'hC7;
        8'hB8: galois_lookup_251 = 8'hB7;
        8'hB9: galois_lookup_251 = 8'h4C;
        8'hBA: galois_lookup_251 = 8'h82;
        8'hBB: galois_lookup_251 = 8'h79;
        8'hBC: galois_lookup_251 = 8'hDD;
        8'hBD: galois_lookup_251 = 8'h26;
        8'hBE: galois_lookup_251 = 8'hE8;
        8'hBF: galois_lookup_251 = 8'h13;
        8'hC0: galois_lookup_251 = 8'hB1;
        8'hC1: galois_lookup_251 = 8'h4A;
        8'hC2: galois_lookup_251 = 8'h84;
        8'hC3: galois_lookup_251 = 8'h7F;
        8'hC4: galois_lookup_251 = 8'hDB;
        8'hC5: galois_lookup_251 = 8'h20;
        8'hC6: galois_lookup_251 = 8'hEE;
        8'hC7: galois_lookup_251 = 8'h15;
        8'hC8: galois_lookup_251 = 8'h65;
        8'hC9: galois_lookup_251 = 8'h9E;
        8'hCA: galois_lookup_251 = 8'h50;
        8'hCB: galois_lookup_251 = 8'hAB;
        8'hCC: galois_lookup_251 = 8'h0F;
        8'hCD: galois_lookup_251 = 8'hF4;
        8'hCE: galois_lookup_251 = 8'h3A;
        8'hCF: galois_lookup_251 = 8'hC1;
        8'hD0: galois_lookup_251 = 8'hDA;
        8'hD1: galois_lookup_251 = 8'h21;
        8'hD2: galois_lookup_251 = 8'hEF;
        8'hD3: galois_lookup_251 = 8'h14;
        8'hD4: galois_lookup_251 = 8'hB0;
        8'hD5: galois_lookup_251 = 8'h4B;
        8'hD6: galois_lookup_251 = 8'h85;
        8'hD7: galois_lookup_251 = 8'h7E;
        8'hD8: galois_lookup_251 = 8'h0E;
        8'hD9: galois_lookup_251 = 8'hF5;
        8'hDA: galois_lookup_251 = 8'h3B;
        8'hDB: galois_lookup_251 = 8'hC0;
        8'hDC: galois_lookup_251 = 8'h64;
        8'hDD: galois_lookup_251 = 8'h9F;
        8'hDE: galois_lookup_251 = 8'h51;
        8'hDF: galois_lookup_251 = 8'hAA;
        8'hE0: galois_lookup_251 = 8'h67;
        8'hE1: galois_lookup_251 = 8'h9C;
        8'hE2: galois_lookup_251 = 8'h52;
        8'hE3: galois_lookup_251 = 8'hA9;
        8'hE4: galois_lookup_251 = 8'h0D;
        8'hE5: galois_lookup_251 = 8'hF6;
        8'hE6: galois_lookup_251 = 8'h38;
        8'hE7: galois_lookup_251 = 8'hC3;
        8'hE8: galois_lookup_251 = 8'hB3;
        8'hE9: galois_lookup_251 = 8'h48;
        8'hEA: galois_lookup_251 = 8'h86;
        8'hEB: galois_lookup_251 = 8'h7D;
        8'hEC: galois_lookup_251 = 8'hD9;
        8'hED: galois_lookup_251 = 8'h22;
        8'hEE: galois_lookup_251 = 8'hEC;
        8'hEF: galois_lookup_251 = 8'h17;
        8'hF0: galois_lookup_251 = 8'h0C;
        8'hF1: galois_lookup_251 = 8'hF7;
        8'hF2: galois_lookup_251 = 8'h39;
        8'hF3: galois_lookup_251 = 8'hC2;
        8'hF4: galois_lookup_251 = 8'h66;
        8'hF5: galois_lookup_251 = 8'h9D;
        8'hF6: galois_lookup_251 = 8'h53;
        8'hF7: galois_lookup_251 = 8'hA8;
        8'hF8: galois_lookup_251 = 8'hD8;
        8'hF9: galois_lookup_251 = 8'h23;
        8'hFA: galois_lookup_251 = 8'hED;
        8'hFB: galois_lookup_251 = 8'h16;
        8'hFC: galois_lookup_251 = 8'hB2;
        8'hFD: galois_lookup_251 = 8'h49;
        8'hFE: galois_lookup_251 = 8'h87;
        8'hFF: galois_lookup_251 = 8'h7C;
    endcase end
endfunction

endmodule
