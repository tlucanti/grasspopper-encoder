`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////
// Company: Miet
// Engineer: Kostya
// 
// Create Date: 19.06.2022 13:19:27
// Design Name: Grasspopper
// Project Name: Grasspopper
// Target Devices: any
// Tool Versions: 2021.1
// Description:
//   header file with lookup tables
//
// Dependencies: None
// 
// Revision: v1.0
//   v0.1 - file Created
//   v1.0 - sbox and galois lookups done
//
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

// `ifndef LOOKUPS_V
// `define LOOKUPS_V

module header();

// // -----------------------------------------------------------------------------
// function automatic [7:0] sbox_lookup;
// /*

// */
//     input   [7:0]   byte;

//     begin case (byte)
//         8'd000: sbox_lookup = 8'hFC;
//         8'd001: sbox_lookup = 8'hEE;
//         8'd002: sbox_lookup = 8'hDD;
//         8'd003: sbox_lookup = 8'h11;
//         8'd004: sbox_lookup = 8'hCF;
//         8'd005: sbox_lookup = 8'h6E;
//         8'd006: sbox_lookup = 8'h31;
//         8'd007: sbox_lookup = 8'h16;
//         8'd008: sbox_lookup = 8'hFB;
//         8'd009: sbox_lookup = 8'hC4;
//         8'd010: sbox_lookup = 8'hFA;
//         8'd011: sbox_lookup = 8'hDA;
//         8'd012: sbox_lookup = 8'h23;
//         8'd013: sbox_lookup = 8'hC5;
//         8'd014: sbox_lookup = 8'h04;
//         8'd015: sbox_lookup = 8'h4D;
//         8'd016: sbox_lookup = 8'hE9;
//         8'd017: sbox_lookup = 8'h77;
//         8'd018: sbox_lookup = 8'hF0;
//         8'd019: sbox_lookup = 8'hDB;
//         8'd020: sbox_lookup = 8'h93;
//         8'd021: sbox_lookup = 8'h2E;
//         8'd022: sbox_lookup = 8'h99;
//         8'd023: sbox_lookup = 8'hBA;
//         8'd024: sbox_lookup = 8'h17;
//         8'd025: sbox_lookup = 8'h36;
//         8'd026: sbox_lookup = 8'hF1;
//         8'd027: sbox_lookup = 8'hBB;
//         8'd028: sbox_lookup = 8'h14;
//         8'd029: sbox_lookup = 8'hCD;
//         8'd030: sbox_lookup = 8'h5F;
//         8'd031: sbox_lookup = 8'hC1;
//         8'd032: sbox_lookup = 8'hF9;
//         8'd033: sbox_lookup = 8'h18;
//         8'd034: sbox_lookup = 8'h65;
//         8'd035: sbox_lookup = 8'h5A;
//         8'd036: sbox_lookup = 8'hE2;
//         8'd037: sbox_lookup = 8'h5C;
//         8'd038: sbox_lookup = 8'hEF;
//         8'd039: sbox_lookup = 8'h21;
//         8'd040: sbox_lookup = 8'h81;
//         8'd041: sbox_lookup = 8'h1C;
//         8'd042: sbox_lookup = 8'h3C;
//         8'd043: sbox_lookup = 8'h42;
//         8'd044: sbox_lookup = 8'h8B;
//         8'd045: sbox_lookup = 8'h01;
//         8'd046: sbox_lookup = 8'h8E;
//         8'd047: sbox_lookup = 8'h4F;
//         8'd048: sbox_lookup = 8'h05;
//         8'd049: sbox_lookup = 8'h84;
//         8'd050: sbox_lookup = 8'h02;
//         8'd051: sbox_lookup = 8'hAE;
//         8'd052: sbox_lookup = 8'hE3;
//         8'd053: sbox_lookup = 8'h6A;
//         8'd054: sbox_lookup = 8'h8F;
//         8'd055: sbox_lookup = 8'hA0;
//         8'd056: sbox_lookup = 8'h06;
//         8'd057: sbox_lookup = 8'h0B;
//         8'd058: sbox_lookup = 8'hED;
//         8'd059: sbox_lookup = 8'h98;
//         8'd060: sbox_lookup = 8'h7F;
//         8'd061: sbox_lookup = 8'hD4;
//         8'd062: sbox_lookup = 8'hD3;
//         8'd063: sbox_lookup = 8'h1F;
//         8'd064: sbox_lookup = 8'hEB;
//         8'd065: sbox_lookup = 8'h34;
//         8'd066: sbox_lookup = 8'h2C;
//         8'd067: sbox_lookup = 8'h51;
//         8'd068: sbox_lookup = 8'hEA;
//         8'd069: sbox_lookup = 8'hC8;
//         8'd070: sbox_lookup = 8'h48;
//         8'd071: sbox_lookup = 8'hAB;
//         8'd072: sbox_lookup = 8'hF2;
//         8'd073: sbox_lookup = 8'h2A;
//         8'd074: sbox_lookup = 8'h68;
//         8'd075: sbox_lookup = 8'hA2;
//         8'd076: sbox_lookup = 8'hFD;
//         8'd077: sbox_lookup = 8'h3A;
//         8'd078: sbox_lookup = 8'hCE;
//         8'd079: sbox_lookup = 8'hCC;
//         8'd080: sbox_lookup = 8'hB5;
//         8'd081: sbox_lookup = 8'h70;
//         8'd082: sbox_lookup = 8'h0E;
//         8'd083: sbox_lookup = 8'h56;
//         8'd084: sbox_lookup = 8'h08;
//         8'd085: sbox_lookup = 8'h0C;
//         8'd086: sbox_lookup = 8'h76;
//         8'd087: sbox_lookup = 8'h12;
//         8'd088: sbox_lookup = 8'hBF;
//         8'd089: sbox_lookup = 8'h72;
//         8'd090: sbox_lookup = 8'h13;
//         8'd091: sbox_lookup = 8'h47;
//         8'd092: sbox_lookup = 8'h9C;
//         8'd093: sbox_lookup = 8'hB7;
//         8'd094: sbox_lookup = 8'h5D;
//         8'd095: sbox_lookup = 8'h87;
//         8'd096: sbox_lookup = 8'h15;
//         8'd097: sbox_lookup = 8'hA1;
//         8'd098: sbox_lookup = 8'h96;
//         8'd099: sbox_lookup = 8'h29;
//         8'd100: sbox_lookup = 8'h10;
//         8'd101: sbox_lookup = 8'h7B;
//         8'd102: sbox_lookup = 8'h9A;
//         8'd103: sbox_lookup = 8'hC7;
//         8'd104: sbox_lookup = 8'hF3;
//         8'd105: sbox_lookup = 8'h91;
//         8'd106: sbox_lookup = 8'h78;
//         8'd107: sbox_lookup = 8'h6F;
//         8'd108: sbox_lookup = 8'h9D;
//         8'd109: sbox_lookup = 8'h9E;
//         8'd110: sbox_lookup = 8'hB2;
//         8'd111: sbox_lookup = 8'hB1;
//         8'd112: sbox_lookup = 8'h32;
//         8'd113: sbox_lookup = 8'h75;
//         8'd114: sbox_lookup = 8'h19;
//         8'd115: sbox_lookup = 8'h3D;
//         8'd116: sbox_lookup = 8'hFF;
//         8'd117: sbox_lookup = 8'h35;
//         8'd118: sbox_lookup = 8'h8A;
//         8'd119: sbox_lookup = 8'h7E;
//         8'd120: sbox_lookup = 8'h6D;
//         8'd121: sbox_lookup = 8'h54;
//         8'd122: sbox_lookup = 8'hC6;
//         8'd123: sbox_lookup = 8'h80;
//         8'd124: sbox_lookup = 8'hC3;
//         8'd125: sbox_lookup = 8'hBD;
//         8'd126: sbox_lookup = 8'h0D;
//         8'd127: sbox_lookup = 8'h57;
//         8'd128: sbox_lookup = 8'hDF;
//         8'd129: sbox_lookup = 8'hF5;
//         8'd130: sbox_lookup = 8'h24;
//         8'd131: sbox_lookup = 8'hA9;
//         8'd132: sbox_lookup = 8'h3E;
//         8'd133: sbox_lookup = 8'hA8;
//         8'd134: sbox_lookup = 8'h43;
//         8'd135: sbox_lookup = 8'hC9;
//         8'd136: sbox_lookup = 8'hD7;
//         8'd137: sbox_lookup = 8'h79;
//         8'd138: sbox_lookup = 8'hD6;
//         8'd139: sbox_lookup = 8'hF6;
//         8'd140: sbox_lookup = 8'h7C;
//         8'd141: sbox_lookup = 8'h22;
//         8'd142: sbox_lookup = 8'hB9;
//         8'd143: sbox_lookup = 8'h03;
//         8'd144: sbox_lookup = 8'hE0;
//         8'd145: sbox_lookup = 8'h0F;
//         8'd146: sbox_lookup = 8'hEC;
//         8'd147: sbox_lookup = 8'hDE;
//         8'd148: sbox_lookup = 8'h7A;
//         8'd149: sbox_lookup = 8'h94;
//         8'd150: sbox_lookup = 8'hB0;
//         8'd151: sbox_lookup = 8'hBC;
//         8'd152: sbox_lookup = 8'hDC;
//         8'd153: sbox_lookup = 8'hE8;
//         8'd154: sbox_lookup = 8'h28;
//         8'd155: sbox_lookup = 8'h50;
//         8'd156: sbox_lookup = 8'h4E;
//         8'd157: sbox_lookup = 8'h33;
//         8'd158: sbox_lookup = 8'h0A;
//         8'd159: sbox_lookup = 8'h4A;
//         8'd160: sbox_lookup = 8'hA7;
//         8'd161: sbox_lookup = 8'h97;
//         8'd162: sbox_lookup = 8'h60;
//         8'd163: sbox_lookup = 8'h73;
//         8'd164: sbox_lookup = 8'h1E;
//         8'd165: sbox_lookup = 8'h00;
//         8'd166: sbox_lookup = 8'h62;
//         8'd167: sbox_lookup = 8'h44;
//         8'd168: sbox_lookup = 8'h1A;
//         8'd169: sbox_lookup = 8'hB8;
//         8'd170: sbox_lookup = 8'h38;
//         8'd171: sbox_lookup = 8'h82;
//         8'd172: sbox_lookup = 8'h64;
//         8'd173: sbox_lookup = 8'h9F;
//         8'd174: sbox_lookup = 8'h26;
//         8'd175: sbox_lookup = 8'h41;
//         8'd176: sbox_lookup = 8'hAD;
//         8'd177: sbox_lookup = 8'h45;
//         8'd178: sbox_lookup = 8'h46;
//         8'd179: sbox_lookup = 8'h92;
//         8'd180: sbox_lookup = 8'h27;
//         8'd181: sbox_lookup = 8'h5E;
//         8'd182: sbox_lookup = 8'h55;
//         8'd183: sbox_lookup = 8'h2F;
//         8'd184: sbox_lookup = 8'h8C;
//         8'd185: sbox_lookup = 8'hA3;
//         8'd186: sbox_lookup = 8'hA5;
//         8'd187: sbox_lookup = 8'h7D;
//         8'd188: sbox_lookup = 8'h69;
//         8'd189: sbox_lookup = 8'hD5;
//         8'd190: sbox_lookup = 8'h95;
//         8'd191: sbox_lookup = 8'h3B;
//         8'd192: sbox_lookup = 8'h07;
//         8'd193: sbox_lookup = 8'h58;
//         8'd194: sbox_lookup = 8'hB3;
//         8'd195: sbox_lookup = 8'h40;
//         8'd196: sbox_lookup = 8'h86;
//         8'd197: sbox_lookup = 8'hAC;
//         8'd198: sbox_lookup = 8'h1D;
//         8'd199: sbox_lookup = 8'hF7;
//         8'd200: sbox_lookup = 8'h30;
//         8'd201: sbox_lookup = 8'h37;
//         8'd202: sbox_lookup = 8'h6B;
//         8'd203: sbox_lookup = 8'hE4;
//         8'd204: sbox_lookup = 8'h88;
//         8'd205: sbox_lookup = 8'hD9;
//         8'd206: sbox_lookup = 8'hE7;
//         8'd207: sbox_lookup = 8'h89;
//         8'd208: sbox_lookup = 8'hE1;
//         8'd209: sbox_lookup = 8'h1B;
//         8'd210: sbox_lookup = 8'h83;
//         8'd211: sbox_lookup = 8'h49;
//         8'd212: sbox_lookup = 8'h4C;
//         8'd213: sbox_lookup = 8'h3F;
//         8'd214: sbox_lookup = 8'hF8;
//         8'd215: sbox_lookup = 8'hFE;
//         8'd216: sbox_lookup = 8'h8D;
//         8'd217: sbox_lookup = 8'h53;
//         8'd218: sbox_lookup = 8'hAA;
//         8'd219: sbox_lookup = 8'h90;
//         8'd220: sbox_lookup = 8'hCA;
//         8'd221: sbox_lookup = 8'hD8;
//         8'd222: sbox_lookup = 8'h85;
//         8'd223: sbox_lookup = 8'h61;
//         8'd224: sbox_lookup = 8'h20;
//         8'd225: sbox_lookup = 8'h71;
//         8'd226: sbox_lookup = 8'h67;
//         8'd227: sbox_lookup = 8'hA4;
//         8'd228: sbox_lookup = 8'h2D;
//         8'd229: sbox_lookup = 8'h2B;
//         8'd230: sbox_lookup = 8'h09;
//         8'd231: sbox_lookup = 8'h5B;
//         8'd232: sbox_lookup = 8'hCB;
//         8'd233: sbox_lookup = 8'h9B;
//         8'd234: sbox_lookup = 8'h25;
//         8'd235: sbox_lookup = 8'hD0;
//         8'd236: sbox_lookup = 8'hBE;
//         8'd237: sbox_lookup = 8'hE5;
//         8'd238: sbox_lookup = 8'h6C;
//         8'd239: sbox_lookup = 8'h52;
//         8'd240: sbox_lookup = 8'h59;
//         8'd241: sbox_lookup = 8'hA6;
//         8'd242: sbox_lookup = 8'h74;
//         8'd243: sbox_lookup = 8'hD2;
//         8'd244: sbox_lookup = 8'hE6;
//         8'd245: sbox_lookup = 8'hF4;
//         8'd246: sbox_lookup = 8'hB4;
//         8'd247: sbox_lookup = 8'hC0;
//         8'd248: sbox_lookup = 8'hD1;
//         8'd249: sbox_lookup = 8'h66;
//         8'd250: sbox_lookup = 8'hAF;
//         8'd251: sbox_lookup = 8'hC2;
//         8'd252: sbox_lookup = 8'h39;
//         8'd253: sbox_lookup = 8'h4B;
//         8'd254: sbox_lookup = 8'h63;
//         8'd255: sbox_lookup = 8'hB6;
//     endcase end
// endfunction

// -----------------------------------------------------------------------------
function automatic [7:0] galois_lookup_016;
/*

*/
    input   [7:0]   byte;

    begin case (byte)
        8'd000: galois_lookup_016 = 8'h00;
        8'd001: galois_lookup_016 = 8'h10;
        8'd002: galois_lookup_016 = 8'h20;
        8'd003: galois_lookup_016 = 8'h30;
        8'd004: galois_lookup_016 = 8'h40;
        8'd005: galois_lookup_016 = 8'h50;
        8'd006: galois_lookup_016 = 8'h60;
        8'd007: galois_lookup_016 = 8'h70;
        8'd008: galois_lookup_016 = 8'h80;
        8'd009: galois_lookup_016 = 8'h90;
        8'd010: galois_lookup_016 = 8'hA0;
        8'd011: galois_lookup_016 = 8'hB0;
        8'd012: galois_lookup_016 = 8'hC0;
        8'd013: galois_lookup_016 = 8'hD0;
        8'd014: galois_lookup_016 = 8'hE0;
        8'd015: galois_lookup_016 = 8'hF0;
        8'd016: galois_lookup_016 = 8'hC3;
        8'd017: galois_lookup_016 = 8'hD3;
        8'd018: galois_lookup_016 = 8'hE3;
        8'd019: galois_lookup_016 = 8'hF3;
        8'd020: galois_lookup_016 = 8'h83;
        8'd021: galois_lookup_016 = 8'h93;
        8'd022: galois_lookup_016 = 8'hA3;
        8'd023: galois_lookup_016 = 8'hB3;
        8'd024: galois_lookup_016 = 8'h43;
        8'd025: galois_lookup_016 = 8'h53;
        8'd026: galois_lookup_016 = 8'h63;
        8'd027: galois_lookup_016 = 8'h73;
        8'd028: galois_lookup_016 = 8'h03;
        8'd029: galois_lookup_016 = 8'h13;
        8'd030: galois_lookup_016 = 8'h23;
        8'd031: galois_lookup_016 = 8'h33;
        8'd032: galois_lookup_016 = 8'h45;
        8'd033: galois_lookup_016 = 8'h55;
        8'd034: galois_lookup_016 = 8'h65;
        8'd035: galois_lookup_016 = 8'h75;
        8'd036: galois_lookup_016 = 8'h05;
        8'd037: galois_lookup_016 = 8'h15;
        8'd038: galois_lookup_016 = 8'h25;
        8'd039: galois_lookup_016 = 8'h35;
        8'd040: galois_lookup_016 = 8'hC5;
        8'd041: galois_lookup_016 = 8'hD5;
        8'd042: galois_lookup_016 = 8'hE5;
        8'd043: galois_lookup_016 = 8'hF5;
        8'd044: galois_lookup_016 = 8'h85;
        8'd045: galois_lookup_016 = 8'h95;
        8'd046: galois_lookup_016 = 8'hA5;
        8'd047: galois_lookup_016 = 8'hB5;
        8'd048: galois_lookup_016 = 8'h86;
        8'd049: galois_lookup_016 = 8'h96;
        8'd050: galois_lookup_016 = 8'hA6;
        8'd051: galois_lookup_016 = 8'hB6;
        8'd052: galois_lookup_016 = 8'hC6;
        8'd053: galois_lookup_016 = 8'hD6;
        8'd054: galois_lookup_016 = 8'hE6;
        8'd055: galois_lookup_016 = 8'hF6;
        8'd056: galois_lookup_016 = 8'h06;
        8'd057: galois_lookup_016 = 8'h16;
        8'd058: galois_lookup_016 = 8'h26;
        8'd059: galois_lookup_016 = 8'h36;
        8'd060: galois_lookup_016 = 8'h46;
        8'd061: galois_lookup_016 = 8'h56;
        8'd062: galois_lookup_016 = 8'h66;
        8'd063: galois_lookup_016 = 8'h76;
        8'd064: galois_lookup_016 = 8'h8A;
        8'd065: galois_lookup_016 = 8'h9A;
        8'd066: galois_lookup_016 = 8'hAA;
        8'd067: galois_lookup_016 = 8'hBA;
        8'd068: galois_lookup_016 = 8'hCA;
        8'd069: galois_lookup_016 = 8'hDA;
        8'd070: galois_lookup_016 = 8'hEA;
        8'd071: galois_lookup_016 = 8'hFA;
        8'd072: galois_lookup_016 = 8'h0A;
        8'd073: galois_lookup_016 = 8'h1A;
        8'd074: galois_lookup_016 = 8'h2A;
        8'd075: galois_lookup_016 = 8'h3A;
        8'd076: galois_lookup_016 = 8'h4A;
        8'd077: galois_lookup_016 = 8'h5A;
        8'd078: galois_lookup_016 = 8'h6A;
        8'd079: galois_lookup_016 = 8'h7A;
        8'd080: galois_lookup_016 = 8'h49;
        8'd081: galois_lookup_016 = 8'h59;
        8'd082: galois_lookup_016 = 8'h69;
        8'd083: galois_lookup_016 = 8'h79;
        8'd084: galois_lookup_016 = 8'h09;
        8'd085: galois_lookup_016 = 8'h19;
        8'd086: galois_lookup_016 = 8'h29;
        8'd087: galois_lookup_016 = 8'h39;
        8'd088: galois_lookup_016 = 8'hC9;
        8'd089: galois_lookup_016 = 8'hD9;
        8'd090: galois_lookup_016 = 8'hE9;
        8'd091: galois_lookup_016 = 8'hF9;
        8'd092: galois_lookup_016 = 8'h89;
        8'd093: galois_lookup_016 = 8'h99;
        8'd094: galois_lookup_016 = 8'hA9;
        8'd095: galois_lookup_016 = 8'hB9;
        8'd096: galois_lookup_016 = 8'hCF;
        8'd097: galois_lookup_016 = 8'hDF;
        8'd098: galois_lookup_016 = 8'hEF;
        8'd099: galois_lookup_016 = 8'hFF;
        8'd100: galois_lookup_016 = 8'h8F;
        8'd101: galois_lookup_016 = 8'h9F;
        8'd102: galois_lookup_016 = 8'hAF;
        8'd103: galois_lookup_016 = 8'hBF;
        8'd104: galois_lookup_016 = 8'h4F;
        8'd105: galois_lookup_016 = 8'h5F;
        8'd106: galois_lookup_016 = 8'h6F;
        8'd107: galois_lookup_016 = 8'h7F;
        8'd108: galois_lookup_016 = 8'h0F;
        8'd109: galois_lookup_016 = 8'h1F;
        8'd110: galois_lookup_016 = 8'h2F;
        8'd111: galois_lookup_016 = 8'h3F;
        8'd112: galois_lookup_016 = 8'h0C;
        8'd113: galois_lookup_016 = 8'h1C;
        8'd114: galois_lookup_016 = 8'h2C;
        8'd115: galois_lookup_016 = 8'h3C;
        8'd116: galois_lookup_016 = 8'h4C;
        8'd117: galois_lookup_016 = 8'h5C;
        8'd118: galois_lookup_016 = 8'h6C;
        8'd119: galois_lookup_016 = 8'h7C;
        8'd120: galois_lookup_016 = 8'h8C;
        8'd121: galois_lookup_016 = 8'h9C;
        8'd122: galois_lookup_016 = 8'hAC;
        8'd123: galois_lookup_016 = 8'hBC;
        8'd124: galois_lookup_016 = 8'hCC;
        8'd125: galois_lookup_016 = 8'hDC;
        8'd126: galois_lookup_016 = 8'hEC;
        8'd127: galois_lookup_016 = 8'hFC;
        8'd128: galois_lookup_016 = 8'hD7;
        8'd129: galois_lookup_016 = 8'hC7;
        8'd130: galois_lookup_016 = 8'hF7;
        8'd131: galois_lookup_016 = 8'hE7;
        8'd132: galois_lookup_016 = 8'h97;
        8'd133: galois_lookup_016 = 8'h87;
        8'd134: galois_lookup_016 = 8'hB7;
        8'd135: galois_lookup_016 = 8'hA7;
        8'd136: galois_lookup_016 = 8'h57;
        8'd137: galois_lookup_016 = 8'h47;
        8'd138: galois_lookup_016 = 8'h77;
        8'd139: galois_lookup_016 = 8'h67;
        8'd140: galois_lookup_016 = 8'h17;
        8'd141: galois_lookup_016 = 8'h07;
        8'd142: galois_lookup_016 = 8'h37;
        8'd143: galois_lookup_016 = 8'h27;
        8'd144: galois_lookup_016 = 8'h14;
        8'd145: galois_lookup_016 = 8'h04;
        8'd146: galois_lookup_016 = 8'h34;
        8'd147: galois_lookup_016 = 8'h24;
        8'd148: galois_lookup_016 = 8'h54;
        8'd149: galois_lookup_016 = 8'h44;
        8'd150: galois_lookup_016 = 8'h74;
        8'd151: galois_lookup_016 = 8'h64;
        8'd152: galois_lookup_016 = 8'h94;
        8'd153: galois_lookup_016 = 8'h84;
        8'd154: galois_lookup_016 = 8'hB4;
        8'd155: galois_lookup_016 = 8'hA4;
        8'd156: galois_lookup_016 = 8'hD4;
        8'd157: galois_lookup_016 = 8'hC4;
        8'd158: galois_lookup_016 = 8'hF4;
        8'd159: galois_lookup_016 = 8'hE4;
        8'd160: galois_lookup_016 = 8'h92;
        8'd161: galois_lookup_016 = 8'h82;
        8'd162: galois_lookup_016 = 8'hB2;
        8'd163: galois_lookup_016 = 8'hA2;
        8'd164: galois_lookup_016 = 8'hD2;
        8'd165: galois_lookup_016 = 8'hC2;
        8'd166: galois_lookup_016 = 8'hF2;
        8'd167: galois_lookup_016 = 8'hE2;
        8'd168: galois_lookup_016 = 8'h12;
        8'd169: galois_lookup_016 = 8'h02;
        8'd170: galois_lookup_016 = 8'h32;
        8'd171: galois_lookup_016 = 8'h22;
        8'd172: galois_lookup_016 = 8'h52;
        8'd173: galois_lookup_016 = 8'h42;
        8'd174: galois_lookup_016 = 8'h72;
        8'd175: galois_lookup_016 = 8'h62;
        8'd176: galois_lookup_016 = 8'h51;
        8'd177: galois_lookup_016 = 8'h41;
        8'd178: galois_lookup_016 = 8'h71;
        8'd179: galois_lookup_016 = 8'h61;
        8'd180: galois_lookup_016 = 8'h11;
        8'd181: galois_lookup_016 = 8'h01;
        8'd182: galois_lookup_016 = 8'h31;
        8'd183: galois_lookup_016 = 8'h21;
        8'd184: galois_lookup_016 = 8'hD1;
        8'd185: galois_lookup_016 = 8'hC1;
        8'd186: galois_lookup_016 = 8'hF1;
        8'd187: galois_lookup_016 = 8'hE1;
        8'd188: galois_lookup_016 = 8'h91;
        8'd189: galois_lookup_016 = 8'h81;
        8'd190: galois_lookup_016 = 8'hB1;
        8'd191: galois_lookup_016 = 8'hA1;
        8'd192: galois_lookup_016 = 8'h5D;
        8'd193: galois_lookup_016 = 8'h4D;
        8'd194: galois_lookup_016 = 8'h7D;
        8'd195: galois_lookup_016 = 8'h6D;
        8'd196: galois_lookup_016 = 8'h1D;
        8'd197: galois_lookup_016 = 8'h0D;
        8'd198: galois_lookup_016 = 8'h3D;
        8'd199: galois_lookup_016 = 8'h2D;
        8'd200: galois_lookup_016 = 8'hDD;
        8'd201: galois_lookup_016 = 8'hCD;
        8'd202: galois_lookup_016 = 8'hFD;
        8'd203: galois_lookup_016 = 8'hED;
        8'd204: galois_lookup_016 = 8'h9D;
        8'd205: galois_lookup_016 = 8'h8D;
        8'd206: galois_lookup_016 = 8'hBD;
        8'd207: galois_lookup_016 = 8'hAD;
        8'd208: galois_lookup_016 = 8'h9E;
        8'd209: galois_lookup_016 = 8'h8E;
        8'd210: galois_lookup_016 = 8'hBE;
        8'd211: galois_lookup_016 = 8'hAE;
        8'd212: galois_lookup_016 = 8'hDE;
        8'd213: galois_lookup_016 = 8'hCE;
        8'd214: galois_lookup_016 = 8'hFE;
        8'd215: galois_lookup_016 = 8'hEE;
        8'd216: galois_lookup_016 = 8'h1E;
        8'd217: galois_lookup_016 = 8'h0E;
        8'd218: galois_lookup_016 = 8'h3E;
        8'd219: galois_lookup_016 = 8'h2E;
        8'd220: galois_lookup_016 = 8'h5E;
        8'd221: galois_lookup_016 = 8'h4E;
        8'd222: galois_lookup_016 = 8'h7E;
        8'd223: galois_lookup_016 = 8'h6E;
        8'd224: galois_lookup_016 = 8'h18;
        8'd225: galois_lookup_016 = 8'h08;
        8'd226: galois_lookup_016 = 8'h38;
        8'd227: galois_lookup_016 = 8'h28;
        8'd228: galois_lookup_016 = 8'h58;
        8'd229: galois_lookup_016 = 8'h48;
        8'd230: galois_lookup_016 = 8'h78;
        8'd231: galois_lookup_016 = 8'h68;
        8'd232: galois_lookup_016 = 8'h98;
        8'd233: galois_lookup_016 = 8'h88;
        8'd234: galois_lookup_016 = 8'hB8;
        8'd235: galois_lookup_016 = 8'hA8;
        8'd236: galois_lookup_016 = 8'hD8;
        8'd237: galois_lookup_016 = 8'hC8;
        8'd238: galois_lookup_016 = 8'hF8;
        8'd239: galois_lookup_016 = 8'hE8;
        8'd240: galois_lookup_016 = 8'hDB;
        8'd241: galois_lookup_016 = 8'hCB;
        8'd242: galois_lookup_016 = 8'hFB;
        8'd243: galois_lookup_016 = 8'hEB;
        8'd244: galois_lookup_016 = 8'h9B;
        8'd245: galois_lookup_016 = 8'h8B;
        8'd246: galois_lookup_016 = 8'hBB;
        8'd247: galois_lookup_016 = 8'hAB;
        8'd248: galois_lookup_016 = 8'h5B;
        8'd249: galois_lookup_016 = 8'h4B;
        8'd250: galois_lookup_016 = 8'h7B;
        8'd251: galois_lookup_016 = 8'h6B;
        8'd252: galois_lookup_016 = 8'h1B;
        8'd253: galois_lookup_016 = 8'h0B;
        8'd254: galois_lookup_016 = 8'h3B;
        8'd255: galois_lookup_016 = 8'h2B;
    endcase end
endfunction

// -----------------------------------------------------------------------------
function automatic [7:0] galois_lookup_032;
/*

*/
    input   [7:0]   byte;

    begin case (byte)
        8'd000: galois_lookup_032 = 8'h00;
        8'd001: galois_lookup_032 = 8'h20;
        8'd002: galois_lookup_032 = 8'h40;
        8'd003: galois_lookup_032 = 8'h60;
        8'd004: galois_lookup_032 = 8'h80;
        8'd005: galois_lookup_032 = 8'hA0;
        8'd006: galois_lookup_032 = 8'hC0;
        8'd007: galois_lookup_032 = 8'hE0;
        8'd008: galois_lookup_032 = 8'hC3;
        8'd009: galois_lookup_032 = 8'hE3;
        8'd010: galois_lookup_032 = 8'h83;
        8'd011: galois_lookup_032 = 8'hA3;
        8'd012: galois_lookup_032 = 8'h43;
        8'd013: galois_lookup_032 = 8'h63;
        8'd014: galois_lookup_032 = 8'h03;
        8'd015: galois_lookup_032 = 8'h23;
        8'd016: galois_lookup_032 = 8'h45;
        8'd017: galois_lookup_032 = 8'h65;
        8'd018: galois_lookup_032 = 8'h05;
        8'd019: galois_lookup_032 = 8'h25;
        8'd020: galois_lookup_032 = 8'hC5;
        8'd021: galois_lookup_032 = 8'hE5;
        8'd022: galois_lookup_032 = 8'h85;
        8'd023: galois_lookup_032 = 8'hA5;
        8'd024: galois_lookup_032 = 8'h86;
        8'd025: galois_lookup_032 = 8'hA6;
        8'd026: galois_lookup_032 = 8'hC6;
        8'd027: galois_lookup_032 = 8'hE6;
        8'd028: galois_lookup_032 = 8'h06;
        8'd029: galois_lookup_032 = 8'h26;
        8'd030: galois_lookup_032 = 8'h46;
        8'd031: galois_lookup_032 = 8'h66;
        8'd032: galois_lookup_032 = 8'h8A;
        8'd033: galois_lookup_032 = 8'hAA;
        8'd034: galois_lookup_032 = 8'hCA;
        8'd035: galois_lookup_032 = 8'hEA;
        8'd036: galois_lookup_032 = 8'h0A;
        8'd037: galois_lookup_032 = 8'h2A;
        8'd038: galois_lookup_032 = 8'h4A;
        8'd039: galois_lookup_032 = 8'h6A;
        8'd040: galois_lookup_032 = 8'h49;
        8'd041: galois_lookup_032 = 8'h69;
        8'd042: galois_lookup_032 = 8'h09;
        8'd043: galois_lookup_032 = 8'h29;
        8'd044: galois_lookup_032 = 8'hC9;
        8'd045: galois_lookup_032 = 8'hE9;
        8'd046: galois_lookup_032 = 8'h89;
        8'd047: galois_lookup_032 = 8'hA9;
        8'd048: galois_lookup_032 = 8'hCF;
        8'd049: galois_lookup_032 = 8'hEF;
        8'd050: galois_lookup_032 = 8'h8F;
        8'd051: galois_lookup_032 = 8'hAF;
        8'd052: galois_lookup_032 = 8'h4F;
        8'd053: galois_lookup_032 = 8'h6F;
        8'd054: galois_lookup_032 = 8'h0F;
        8'd055: galois_lookup_032 = 8'h2F;
        8'd056: galois_lookup_032 = 8'h0C;
        8'd057: galois_lookup_032 = 8'h2C;
        8'd058: galois_lookup_032 = 8'h4C;
        8'd059: galois_lookup_032 = 8'h6C;
        8'd060: galois_lookup_032 = 8'h8C;
        8'd061: galois_lookup_032 = 8'hAC;
        8'd062: galois_lookup_032 = 8'hCC;
        8'd063: galois_lookup_032 = 8'hEC;
        8'd064: galois_lookup_032 = 8'hD7;
        8'd065: galois_lookup_032 = 8'hF7;
        8'd066: galois_lookup_032 = 8'h97;
        8'd067: galois_lookup_032 = 8'hB7;
        8'd068: galois_lookup_032 = 8'h57;
        8'd069: galois_lookup_032 = 8'h77;
        8'd070: galois_lookup_032 = 8'h17;
        8'd071: galois_lookup_032 = 8'h37;
        8'd072: galois_lookup_032 = 8'h14;
        8'd073: galois_lookup_032 = 8'h34;
        8'd074: galois_lookup_032 = 8'h54;
        8'd075: galois_lookup_032 = 8'h74;
        8'd076: galois_lookup_032 = 8'h94;
        8'd077: galois_lookup_032 = 8'hB4;
        8'd078: galois_lookup_032 = 8'hD4;
        8'd079: galois_lookup_032 = 8'hF4;
        8'd080: galois_lookup_032 = 8'h92;
        8'd081: galois_lookup_032 = 8'hB2;
        8'd082: galois_lookup_032 = 8'hD2;
        8'd083: galois_lookup_032 = 8'hF2;
        8'd084: galois_lookup_032 = 8'h12;
        8'd085: galois_lookup_032 = 8'h32;
        8'd086: galois_lookup_032 = 8'h52;
        8'd087: galois_lookup_032 = 8'h72;
        8'd088: galois_lookup_032 = 8'h51;
        8'd089: galois_lookup_032 = 8'h71;
        8'd090: galois_lookup_032 = 8'h11;
        8'd091: galois_lookup_032 = 8'h31;
        8'd092: galois_lookup_032 = 8'hD1;
        8'd093: galois_lookup_032 = 8'hF1;
        8'd094: galois_lookup_032 = 8'h91;
        8'd095: galois_lookup_032 = 8'hB1;
        8'd096: galois_lookup_032 = 8'h5D;
        8'd097: galois_lookup_032 = 8'h7D;
        8'd098: galois_lookup_032 = 8'h1D;
        8'd099: galois_lookup_032 = 8'h3D;
        8'd100: galois_lookup_032 = 8'hDD;
        8'd101: galois_lookup_032 = 8'hFD;
        8'd102: galois_lookup_032 = 8'h9D;
        8'd103: galois_lookup_032 = 8'hBD;
        8'd104: galois_lookup_032 = 8'h9E;
        8'd105: galois_lookup_032 = 8'hBE;
        8'd106: galois_lookup_032 = 8'hDE;
        8'd107: galois_lookup_032 = 8'hFE;
        8'd108: galois_lookup_032 = 8'h1E;
        8'd109: galois_lookup_032 = 8'h3E;
        8'd110: galois_lookup_032 = 8'h5E;
        8'd111: galois_lookup_032 = 8'h7E;
        8'd112: galois_lookup_032 = 8'h18;
        8'd113: galois_lookup_032 = 8'h38;
        8'd114: galois_lookup_032 = 8'h58;
        8'd115: galois_lookup_032 = 8'h78;
        8'd116: galois_lookup_032 = 8'h98;
        8'd117: galois_lookup_032 = 8'hB8;
        8'd118: galois_lookup_032 = 8'hD8;
        8'd119: galois_lookup_032 = 8'hF8;
        8'd120: galois_lookup_032 = 8'hDB;
        8'd121: galois_lookup_032 = 8'hFB;
        8'd122: galois_lookup_032 = 8'h9B;
        8'd123: galois_lookup_032 = 8'hBB;
        8'd124: galois_lookup_032 = 8'h5B;
        8'd125: galois_lookup_032 = 8'h7B;
        8'd126: galois_lookup_032 = 8'h1B;
        8'd127: galois_lookup_032 = 8'h3B;
        8'd128: galois_lookup_032 = 8'h6D;
        8'd129: galois_lookup_032 = 8'h4D;
        8'd130: galois_lookup_032 = 8'h2D;
        8'd131: galois_lookup_032 = 8'h0D;
        8'd132: galois_lookup_032 = 8'hED;
        8'd133: galois_lookup_032 = 8'hCD;
        8'd134: galois_lookup_032 = 8'hAD;
        8'd135: galois_lookup_032 = 8'h8D;
        8'd136: galois_lookup_032 = 8'hAE;
        8'd137: galois_lookup_032 = 8'h8E;
        8'd138: galois_lookup_032 = 8'hEE;
        8'd139: galois_lookup_032 = 8'hCE;
        8'd140: galois_lookup_032 = 8'h2E;
        8'd141: galois_lookup_032 = 8'h0E;
        8'd142: galois_lookup_032 = 8'h6E;
        8'd143: galois_lookup_032 = 8'h4E;
        8'd144: galois_lookup_032 = 8'h28;
        8'd145: galois_lookup_032 = 8'h08;
        8'd146: galois_lookup_032 = 8'h68;
        8'd147: galois_lookup_032 = 8'h48;
        8'd148: galois_lookup_032 = 8'hA8;
        8'd149: galois_lookup_032 = 8'h88;
        8'd150: galois_lookup_032 = 8'hE8;
        8'd151: galois_lookup_032 = 8'hC8;
        8'd152: galois_lookup_032 = 8'hEB;
        8'd153: galois_lookup_032 = 8'hCB;
        8'd154: galois_lookup_032 = 8'hAB;
        8'd155: galois_lookup_032 = 8'h8B;
        8'd156: galois_lookup_032 = 8'h6B;
        8'd157: galois_lookup_032 = 8'h4B;
        8'd158: galois_lookup_032 = 8'h2B;
        8'd159: galois_lookup_032 = 8'h0B;
        8'd160: galois_lookup_032 = 8'hE7;
        8'd161: galois_lookup_032 = 8'hC7;
        8'd162: galois_lookup_032 = 8'hA7;
        8'd163: galois_lookup_032 = 8'h87;
        8'd164: galois_lookup_032 = 8'h67;
        8'd165: galois_lookup_032 = 8'h47;
        8'd166: galois_lookup_032 = 8'h27;
        8'd167: galois_lookup_032 = 8'h07;
        8'd168: galois_lookup_032 = 8'h24;
        8'd169: galois_lookup_032 = 8'h04;
        8'd170: galois_lookup_032 = 8'h64;
        8'd171: galois_lookup_032 = 8'h44;
        8'd172: galois_lookup_032 = 8'hA4;
        8'd173: galois_lookup_032 = 8'h84;
        8'd174: galois_lookup_032 = 8'hE4;
        8'd175: galois_lookup_032 = 8'hC4;
        8'd176: galois_lookup_032 = 8'hA2;
        8'd177: galois_lookup_032 = 8'h82;
        8'd178: galois_lookup_032 = 8'hE2;
        8'd179: galois_lookup_032 = 8'hC2;
        8'd180: galois_lookup_032 = 8'h22;
        8'd181: galois_lookup_032 = 8'h02;
        8'd182: galois_lookup_032 = 8'h62;
        8'd183: galois_lookup_032 = 8'h42;
        8'd184: galois_lookup_032 = 8'h61;
        8'd185: galois_lookup_032 = 8'h41;
        8'd186: galois_lookup_032 = 8'h21;
        8'd187: galois_lookup_032 = 8'h01;
        8'd188: galois_lookup_032 = 8'hE1;
        8'd189: galois_lookup_032 = 8'hC1;
        8'd190: galois_lookup_032 = 8'hA1;
        8'd191: galois_lookup_032 = 8'h81;
        8'd192: galois_lookup_032 = 8'hBA;
        8'd193: galois_lookup_032 = 8'h9A;
        8'd194: galois_lookup_032 = 8'hFA;
        8'd195: galois_lookup_032 = 8'hDA;
        8'd196: galois_lookup_032 = 8'h3A;
        8'd197: galois_lookup_032 = 8'h1A;
        8'd198: galois_lookup_032 = 8'h7A;
        8'd199: galois_lookup_032 = 8'h5A;
        8'd200: galois_lookup_032 = 8'h79;
        8'd201: galois_lookup_032 = 8'h59;
        8'd202: galois_lookup_032 = 8'h39;
        8'd203: galois_lookup_032 = 8'h19;
        8'd204: galois_lookup_032 = 8'hF9;
        8'd205: galois_lookup_032 = 8'hD9;
        8'd206: galois_lookup_032 = 8'hB9;
        8'd207: galois_lookup_032 = 8'h99;
        8'd208: galois_lookup_032 = 8'hFF;
        8'd209: galois_lookup_032 = 8'hDF;
        8'd210: galois_lookup_032 = 8'hBF;
        8'd211: galois_lookup_032 = 8'h9F;
        8'd212: galois_lookup_032 = 8'h7F;
        8'd213: galois_lookup_032 = 8'h5F;
        8'd214: galois_lookup_032 = 8'h3F;
        8'd215: galois_lookup_032 = 8'h1F;
        8'd216: galois_lookup_032 = 8'h3C;
        8'd217: galois_lookup_032 = 8'h1C;
        8'd218: galois_lookup_032 = 8'h7C;
        8'd219: galois_lookup_032 = 8'h5C;
        8'd220: galois_lookup_032 = 8'hBC;
        8'd221: galois_lookup_032 = 8'h9C;
        8'd222: galois_lookup_032 = 8'hFC;
        8'd223: galois_lookup_032 = 8'hDC;
        8'd224: galois_lookup_032 = 8'h30;
        8'd225: galois_lookup_032 = 8'h10;
        8'd226: galois_lookup_032 = 8'h70;
        8'd227: galois_lookup_032 = 8'h50;
        8'd228: galois_lookup_032 = 8'hB0;
        8'd229: galois_lookup_032 = 8'h90;
        8'd230: galois_lookup_032 = 8'hF0;
        8'd231: galois_lookup_032 = 8'hD0;
        8'd232: galois_lookup_032 = 8'hF3;
        8'd233: galois_lookup_032 = 8'hD3;
        8'd234: galois_lookup_032 = 8'hB3;
        8'd235: galois_lookup_032 = 8'h93;
        8'd236: galois_lookup_032 = 8'h73;
        8'd237: galois_lookup_032 = 8'h53;
        8'd238: galois_lookup_032 = 8'h33;
        8'd239: galois_lookup_032 = 8'h13;
        8'd240: galois_lookup_032 = 8'h75;
        8'd241: galois_lookup_032 = 8'h55;
        8'd242: galois_lookup_032 = 8'h35;
        8'd243: galois_lookup_032 = 8'h15;
        8'd244: galois_lookup_032 = 8'hF5;
        8'd245: galois_lookup_032 = 8'hD5;
        8'd246: galois_lookup_032 = 8'hB5;
        8'd247: galois_lookup_032 = 8'h95;
        8'd248: galois_lookup_032 = 8'hB6;
        8'd249: galois_lookup_032 = 8'h96;
        8'd250: galois_lookup_032 = 8'hF6;
        8'd251: galois_lookup_032 = 8'hD6;
        8'd252: galois_lookup_032 = 8'h36;
        8'd253: galois_lookup_032 = 8'h16;
        8'd254: galois_lookup_032 = 8'h76;
        8'd255: galois_lookup_032 = 8'h56;
    endcase end
endfunction

// -----------------------------------------------------------------------------
function automatic [7:0] galois_lookup_133;
/*

*/
    input   [7:0]   byte;

    begin case (byte)
        8'd000: galois_lookup_133 = 8'h00;
        8'd001: galois_lookup_133 = 8'h85;
        8'd002: galois_lookup_133 = 8'hC9;
        8'd003: galois_lookup_133 = 8'h4C;
        8'd004: galois_lookup_133 = 8'h51;
        8'd005: galois_lookup_133 = 8'hD4;
        8'd006: galois_lookup_133 = 8'h98;
        8'd007: galois_lookup_133 = 8'h1D;
        8'd008: galois_lookup_133 = 8'hA2;
        8'd009: galois_lookup_133 = 8'h27;
        8'd010: galois_lookup_133 = 8'h6B;
        8'd011: galois_lookup_133 = 8'hEE;
        8'd012: galois_lookup_133 = 8'hF3;
        8'd013: galois_lookup_133 = 8'h76;
        8'd014: galois_lookup_133 = 8'h3A;
        8'd015: galois_lookup_133 = 8'hBF;
        8'd016: galois_lookup_133 = 8'h87;
        8'd017: galois_lookup_133 = 8'h02;
        8'd018: galois_lookup_133 = 8'h4E;
        8'd019: galois_lookup_133 = 8'hCB;
        8'd020: galois_lookup_133 = 8'hD6;
        8'd021: galois_lookup_133 = 8'h53;
        8'd022: galois_lookup_133 = 8'h1F;
        8'd023: galois_lookup_133 = 8'h9A;
        8'd024: galois_lookup_133 = 8'h25;
        8'd025: galois_lookup_133 = 8'hA0;
        8'd026: galois_lookup_133 = 8'hEC;
        8'd027: galois_lookup_133 = 8'h69;
        8'd028: galois_lookup_133 = 8'h74;
        8'd029: galois_lookup_133 = 8'hF1;
        8'd030: galois_lookup_133 = 8'hBD;
        8'd031: galois_lookup_133 = 8'h38;
        8'd032: galois_lookup_133 = 8'hCD;
        8'd033: galois_lookup_133 = 8'h48;
        8'd034: galois_lookup_133 = 8'h04;
        8'd035: galois_lookup_133 = 8'h81;
        8'd036: galois_lookup_133 = 8'h9C;
        8'd037: galois_lookup_133 = 8'h19;
        8'd038: galois_lookup_133 = 8'h55;
        8'd039: galois_lookup_133 = 8'hD0;
        8'd040: galois_lookup_133 = 8'h6F;
        8'd041: galois_lookup_133 = 8'hEA;
        8'd042: galois_lookup_133 = 8'hA6;
        8'd043: galois_lookup_133 = 8'h23;
        8'd044: galois_lookup_133 = 8'h3E;
        8'd045: galois_lookup_133 = 8'hBB;
        8'd046: galois_lookup_133 = 8'hF7;
        8'd047: galois_lookup_133 = 8'h72;
        8'd048: galois_lookup_133 = 8'h4A;
        8'd049: galois_lookup_133 = 8'hCF;
        8'd050: galois_lookup_133 = 8'h83;
        8'd051: galois_lookup_133 = 8'h06;
        8'd052: galois_lookup_133 = 8'h1B;
        8'd053: galois_lookup_133 = 8'h9E;
        8'd054: galois_lookup_133 = 8'hD2;
        8'd055: galois_lookup_133 = 8'h57;
        8'd056: galois_lookup_133 = 8'hE8;
        8'd057: galois_lookup_133 = 8'h6D;
        8'd058: galois_lookup_133 = 8'h21;
        8'd059: galois_lookup_133 = 8'hA4;
        8'd060: galois_lookup_133 = 8'hB9;
        8'd061: galois_lookup_133 = 8'h3C;
        8'd062: galois_lookup_133 = 8'h70;
        8'd063: galois_lookup_133 = 8'hF5;
        8'd064: galois_lookup_133 = 8'h59;
        8'd065: galois_lookup_133 = 8'hDC;
        8'd066: galois_lookup_133 = 8'h90;
        8'd067: galois_lookup_133 = 8'h15;
        8'd068: galois_lookup_133 = 8'h08;
        8'd069: galois_lookup_133 = 8'h8D;
        8'd070: galois_lookup_133 = 8'hC1;
        8'd071: galois_lookup_133 = 8'h44;
        8'd072: galois_lookup_133 = 8'hFB;
        8'd073: galois_lookup_133 = 8'h7E;
        8'd074: galois_lookup_133 = 8'h32;
        8'd075: galois_lookup_133 = 8'hB7;
        8'd076: galois_lookup_133 = 8'hAA;
        8'd077: galois_lookup_133 = 8'h2F;
        8'd078: galois_lookup_133 = 8'h63;
        8'd079: galois_lookup_133 = 8'hE6;
        8'd080: galois_lookup_133 = 8'hDE;
        8'd081: galois_lookup_133 = 8'h5B;
        8'd082: galois_lookup_133 = 8'h17;
        8'd083: galois_lookup_133 = 8'h92;
        8'd084: galois_lookup_133 = 8'h8F;
        8'd085: galois_lookup_133 = 8'h0A;
        8'd086: galois_lookup_133 = 8'h46;
        8'd087: galois_lookup_133 = 8'hC3;
        8'd088: galois_lookup_133 = 8'h7C;
        8'd089: galois_lookup_133 = 8'hF9;
        8'd090: galois_lookup_133 = 8'hB5;
        8'd091: galois_lookup_133 = 8'h30;
        8'd092: galois_lookup_133 = 8'h2D;
        8'd093: galois_lookup_133 = 8'hA8;
        8'd094: galois_lookup_133 = 8'hE4;
        8'd095: galois_lookup_133 = 8'h61;
        8'd096: galois_lookup_133 = 8'h94;
        8'd097: galois_lookup_133 = 8'h11;
        8'd098: galois_lookup_133 = 8'h5D;
        8'd099: galois_lookup_133 = 8'hD8;
        8'd100: galois_lookup_133 = 8'hC5;
        8'd101: galois_lookup_133 = 8'h40;
        8'd102: galois_lookup_133 = 8'h0C;
        8'd103: galois_lookup_133 = 8'h89;
        8'd104: galois_lookup_133 = 8'h36;
        8'd105: galois_lookup_133 = 8'hB3;
        8'd106: galois_lookup_133 = 8'hFF;
        8'd107: galois_lookup_133 = 8'h7A;
        8'd108: galois_lookup_133 = 8'h67;
        8'd109: galois_lookup_133 = 8'hE2;
        8'd110: galois_lookup_133 = 8'hAE;
        8'd111: galois_lookup_133 = 8'h2B;
        8'd112: galois_lookup_133 = 8'h13;
        8'd113: galois_lookup_133 = 8'h96;
        8'd114: galois_lookup_133 = 8'hDA;
        8'd115: galois_lookup_133 = 8'h5F;
        8'd116: galois_lookup_133 = 8'h42;
        8'd117: galois_lookup_133 = 8'hC7;
        8'd118: galois_lookup_133 = 8'h8B;
        8'd119: galois_lookup_133 = 8'h0E;
        8'd120: galois_lookup_133 = 8'hB1;
        8'd121: galois_lookup_133 = 8'h34;
        8'd122: galois_lookup_133 = 8'h78;
        8'd123: galois_lookup_133 = 8'hFD;
        8'd124: galois_lookup_133 = 8'hE0;
        8'd125: galois_lookup_133 = 8'h65;
        8'd126: galois_lookup_133 = 8'h29;
        8'd127: galois_lookup_133 = 8'hAC;
        8'd128: galois_lookup_133 = 8'hB2;
        8'd129: galois_lookup_133 = 8'h37;
        8'd130: galois_lookup_133 = 8'h7B;
        8'd131: galois_lookup_133 = 8'hFE;
        8'd132: galois_lookup_133 = 8'hE3;
        8'd133: galois_lookup_133 = 8'h66;
        8'd134: galois_lookup_133 = 8'h2A;
        8'd135: galois_lookup_133 = 8'hAF;
        8'd136: galois_lookup_133 = 8'h10;
        8'd137: galois_lookup_133 = 8'h95;
        8'd138: galois_lookup_133 = 8'hD9;
        8'd139: galois_lookup_133 = 8'h5C;
        8'd140: galois_lookup_133 = 8'h41;
        8'd141: galois_lookup_133 = 8'hC4;
        8'd142: galois_lookup_133 = 8'h88;
        8'd143: galois_lookup_133 = 8'h0D;
        8'd144: galois_lookup_133 = 8'h35;
        8'd145: galois_lookup_133 = 8'hB0;
        8'd146: galois_lookup_133 = 8'hFC;
        8'd147: galois_lookup_133 = 8'h79;
        8'd148: galois_lookup_133 = 8'h64;
        8'd149: galois_lookup_133 = 8'hE1;
        8'd150: galois_lookup_133 = 8'hAD;
        8'd151: galois_lookup_133 = 8'h28;
        8'd152: galois_lookup_133 = 8'h97;
        8'd153: galois_lookup_133 = 8'h12;
        8'd154: galois_lookup_133 = 8'h5E;
        8'd155: galois_lookup_133 = 8'hDB;
        8'd156: galois_lookup_133 = 8'hC6;
        8'd157: galois_lookup_133 = 8'h43;
        8'd158: galois_lookup_133 = 8'h0F;
        8'd159: galois_lookup_133 = 8'h8A;
        8'd160: galois_lookup_133 = 8'h7F;
        8'd161: galois_lookup_133 = 8'hFA;
        8'd162: galois_lookup_133 = 8'hB6;
        8'd163: galois_lookup_133 = 8'h33;
        8'd164: galois_lookup_133 = 8'h2E;
        8'd165: galois_lookup_133 = 8'hAB;
        8'd166: galois_lookup_133 = 8'hE7;
        8'd167: galois_lookup_133 = 8'h62;
        8'd168: galois_lookup_133 = 8'hDD;
        8'd169: galois_lookup_133 = 8'h58;
        8'd170: galois_lookup_133 = 8'h14;
        8'd171: galois_lookup_133 = 8'h91;
        8'd172: galois_lookup_133 = 8'h8C;
        8'd173: galois_lookup_133 = 8'h09;
        8'd174: galois_lookup_133 = 8'h45;
        8'd175: galois_lookup_133 = 8'hC0;
        8'd176: galois_lookup_133 = 8'hF8;
        8'd177: galois_lookup_133 = 8'h7D;
        8'd178: galois_lookup_133 = 8'h31;
        8'd179: galois_lookup_133 = 8'hB4;
        8'd180: galois_lookup_133 = 8'hA9;
        8'd181: galois_lookup_133 = 8'h2C;
        8'd182: galois_lookup_133 = 8'h60;
        8'd183: galois_lookup_133 = 8'hE5;
        8'd184: galois_lookup_133 = 8'h5A;
        8'd185: galois_lookup_133 = 8'hDF;
        8'd186: galois_lookup_133 = 8'h93;
        8'd187: galois_lookup_133 = 8'h16;
        8'd188: galois_lookup_133 = 8'h0B;
        8'd189: galois_lookup_133 = 8'h8E;
        8'd190: galois_lookup_133 = 8'hC2;
        8'd191: galois_lookup_133 = 8'h47;
        8'd192: galois_lookup_133 = 8'hEB;
        8'd193: galois_lookup_133 = 8'h6E;
        8'd194: galois_lookup_133 = 8'h22;
        8'd195: galois_lookup_133 = 8'hA7;
        8'd196: galois_lookup_133 = 8'hBA;
        8'd197: galois_lookup_133 = 8'h3F;
        8'd198: galois_lookup_133 = 8'h73;
        8'd199: galois_lookup_133 = 8'hF6;
        8'd200: galois_lookup_133 = 8'h49;
        8'd201: galois_lookup_133 = 8'hCC;
        8'd202: galois_lookup_133 = 8'h80;
        8'd203: galois_lookup_133 = 8'h05;
        8'd204: galois_lookup_133 = 8'h18;
        8'd205: galois_lookup_133 = 8'h9D;
        8'd206: galois_lookup_133 = 8'hD1;
        8'd207: galois_lookup_133 = 8'h54;
        8'd208: galois_lookup_133 = 8'h6C;
        8'd209: galois_lookup_133 = 8'hE9;
        8'd210: galois_lookup_133 = 8'hA5;
        8'd211: galois_lookup_133 = 8'h20;
        8'd212: galois_lookup_133 = 8'h3D;
        8'd213: galois_lookup_133 = 8'hB8;
        8'd214: galois_lookup_133 = 8'hF4;
        8'd215: galois_lookup_133 = 8'h71;
        8'd216: galois_lookup_133 = 8'hCE;
        8'd217: galois_lookup_133 = 8'h4B;
        8'd218: galois_lookup_133 = 8'h07;
        8'd219: galois_lookup_133 = 8'h82;
        8'd220: galois_lookup_133 = 8'h9F;
        8'd221: galois_lookup_133 = 8'h1A;
        8'd222: galois_lookup_133 = 8'h56;
        8'd223: galois_lookup_133 = 8'hD3;
        8'd224: galois_lookup_133 = 8'h26;
        8'd225: galois_lookup_133 = 8'hA3;
        8'd226: galois_lookup_133 = 8'hEF;
        8'd227: galois_lookup_133 = 8'h6A;
        8'd228: galois_lookup_133 = 8'h77;
        8'd229: galois_lookup_133 = 8'hF2;
        8'd230: galois_lookup_133 = 8'hBE;
        8'd231: galois_lookup_133 = 8'h3B;
        8'd232: galois_lookup_133 = 8'h84;
        8'd233: galois_lookup_133 = 8'h01;
        8'd234: galois_lookup_133 = 8'h4D;
        8'd235: galois_lookup_133 = 8'hC8;
        8'd236: galois_lookup_133 = 8'hD5;
        8'd237: galois_lookup_133 = 8'h50;
        8'd238: galois_lookup_133 = 8'h1C;
        8'd239: galois_lookup_133 = 8'h99;
        8'd240: galois_lookup_133 = 8'hA1;
        8'd241: galois_lookup_133 = 8'h24;
        8'd242: galois_lookup_133 = 8'h68;
        8'd243: galois_lookup_133 = 8'hED;
        8'd244: galois_lookup_133 = 8'hF0;
        8'd245: galois_lookup_133 = 8'h75;
        8'd246: galois_lookup_133 = 8'h39;
        8'd247: galois_lookup_133 = 8'hBC;
        8'd248: galois_lookup_133 = 8'h03;
        8'd249: galois_lookup_133 = 8'h86;
        8'd250: galois_lookup_133 = 8'hCA;
        8'd251: galois_lookup_133 = 8'h4F;
        8'd252: galois_lookup_133 = 8'h52;
        8'd253: galois_lookup_133 = 8'hD7;
        8'd254: galois_lookup_133 = 8'h9B;
        8'd255: galois_lookup_133 = 8'h1E;
    endcase end
endfunction

// -----------------------------------------------------------------------------
function automatic [7:0] galois_lookup_148;
/*

*/
    input   [7:0]   byte;

    begin case (byte)
        8'd000: galois_lookup_148 = 8'h00;
        8'd001: galois_lookup_148 = 8'h94;
        8'd002: galois_lookup_148 = 8'hEB;
        8'd003: galois_lookup_148 = 8'h7F;
        8'd004: galois_lookup_148 = 8'h15;
        8'd005: galois_lookup_148 = 8'h81;
        8'd006: galois_lookup_148 = 8'hFE;
        8'd007: galois_lookup_148 = 8'h6A;
        8'd008: galois_lookup_148 = 8'h2A;
        8'd009: galois_lookup_148 = 8'hBE;
        8'd010: galois_lookup_148 = 8'hC1;
        8'd011: galois_lookup_148 = 8'h55;
        8'd012: galois_lookup_148 = 8'h3F;
        8'd013: galois_lookup_148 = 8'hAB;
        8'd014: galois_lookup_148 = 8'hD4;
        8'd015: galois_lookup_148 = 8'h40;
        8'd016: galois_lookup_148 = 8'h54;
        8'd017: galois_lookup_148 = 8'hC0;
        8'd018: galois_lookup_148 = 8'hBF;
        8'd019: galois_lookup_148 = 8'h2B;
        8'd020: galois_lookup_148 = 8'h41;
        8'd021: galois_lookup_148 = 8'hD5;
        8'd022: galois_lookup_148 = 8'hAA;
        8'd023: galois_lookup_148 = 8'h3E;
        8'd024: galois_lookup_148 = 8'h7E;
        8'd025: galois_lookup_148 = 8'hEA;
        8'd026: galois_lookup_148 = 8'h95;
        8'd027: galois_lookup_148 = 8'h01;
        8'd028: galois_lookup_148 = 8'h6B;
        8'd029: galois_lookup_148 = 8'hFF;
        8'd030: galois_lookup_148 = 8'h80;
        8'd031: galois_lookup_148 = 8'h14;
        8'd032: galois_lookup_148 = 8'hA8;
        8'd033: galois_lookup_148 = 8'h3C;
        8'd034: galois_lookup_148 = 8'h43;
        8'd035: galois_lookup_148 = 8'hD7;
        8'd036: galois_lookup_148 = 8'hBD;
        8'd037: galois_lookup_148 = 8'h29;
        8'd038: galois_lookup_148 = 8'h56;
        8'd039: galois_lookup_148 = 8'hC2;
        8'd040: galois_lookup_148 = 8'h82;
        8'd041: galois_lookup_148 = 8'h16;
        8'd042: galois_lookup_148 = 8'h69;
        8'd043: galois_lookup_148 = 8'hFD;
        8'd044: galois_lookup_148 = 8'h97;
        8'd045: galois_lookup_148 = 8'h03;
        8'd046: galois_lookup_148 = 8'h7C;
        8'd047: galois_lookup_148 = 8'hE8;
        8'd048: galois_lookup_148 = 8'hFC;
        8'd049: galois_lookup_148 = 8'h68;
        8'd050: galois_lookup_148 = 8'h17;
        8'd051: galois_lookup_148 = 8'h83;
        8'd052: galois_lookup_148 = 8'hE9;
        8'd053: galois_lookup_148 = 8'h7D;
        8'd054: galois_lookup_148 = 8'h02;
        8'd055: galois_lookup_148 = 8'h96;
        8'd056: galois_lookup_148 = 8'hD6;
        8'd057: galois_lookup_148 = 8'h42;
        8'd058: galois_lookup_148 = 8'h3D;
        8'd059: galois_lookup_148 = 8'hA9;
        8'd060: galois_lookup_148 = 8'hC3;
        8'd061: galois_lookup_148 = 8'h57;
        8'd062: galois_lookup_148 = 8'h28;
        8'd063: galois_lookup_148 = 8'hBC;
        8'd064: galois_lookup_148 = 8'h93;
        8'd065: galois_lookup_148 = 8'h07;
        8'd066: galois_lookup_148 = 8'h78;
        8'd067: galois_lookup_148 = 8'hEC;
        8'd068: galois_lookup_148 = 8'h86;
        8'd069: galois_lookup_148 = 8'h12;
        8'd070: galois_lookup_148 = 8'h6D;
        8'd071: galois_lookup_148 = 8'hF9;
        8'd072: galois_lookup_148 = 8'hB9;
        8'd073: galois_lookup_148 = 8'h2D;
        8'd074: galois_lookup_148 = 8'h52;
        8'd075: galois_lookup_148 = 8'hC6;
        8'd076: galois_lookup_148 = 8'hAC;
        8'd077: galois_lookup_148 = 8'h38;
        8'd078: galois_lookup_148 = 8'h47;
        8'd079: galois_lookup_148 = 8'hD3;
        8'd080: galois_lookup_148 = 8'hC7;
        8'd081: galois_lookup_148 = 8'h53;
        8'd082: galois_lookup_148 = 8'h2C;
        8'd083: galois_lookup_148 = 8'hB8;
        8'd084: galois_lookup_148 = 8'hD2;
        8'd085: galois_lookup_148 = 8'h46;
        8'd086: galois_lookup_148 = 8'h39;
        8'd087: galois_lookup_148 = 8'hAD;
        8'd088: galois_lookup_148 = 8'hED;
        8'd089: galois_lookup_148 = 8'h79;
        8'd090: galois_lookup_148 = 8'h06;
        8'd091: galois_lookup_148 = 8'h92;
        8'd092: galois_lookup_148 = 8'hF8;
        8'd093: galois_lookup_148 = 8'h6C;
        8'd094: galois_lookup_148 = 8'h13;
        8'd095: galois_lookup_148 = 8'h87;
        8'd096: galois_lookup_148 = 8'h3B;
        8'd097: galois_lookup_148 = 8'hAF;
        8'd098: galois_lookup_148 = 8'hD0;
        8'd099: galois_lookup_148 = 8'h44;
        8'd100: galois_lookup_148 = 8'h2E;
        8'd101: galois_lookup_148 = 8'hBA;
        8'd102: galois_lookup_148 = 8'hC5;
        8'd103: galois_lookup_148 = 8'h51;
        8'd104: galois_lookup_148 = 8'h11;
        8'd105: galois_lookup_148 = 8'h85;
        8'd106: galois_lookup_148 = 8'hFA;
        8'd107: galois_lookup_148 = 8'h6E;
        8'd108: galois_lookup_148 = 8'h04;
        8'd109: galois_lookup_148 = 8'h90;
        8'd110: galois_lookup_148 = 8'hEF;
        8'd111: galois_lookup_148 = 8'h7B;
        8'd112: galois_lookup_148 = 8'h6F;
        8'd113: galois_lookup_148 = 8'hFB;
        8'd114: galois_lookup_148 = 8'h84;
        8'd115: galois_lookup_148 = 8'h10;
        8'd116: galois_lookup_148 = 8'h7A;
        8'd117: galois_lookup_148 = 8'hEE;
        8'd118: galois_lookup_148 = 8'h91;
        8'd119: galois_lookup_148 = 8'h05;
        8'd120: galois_lookup_148 = 8'h45;
        8'd121: galois_lookup_148 = 8'hD1;
        8'd122: galois_lookup_148 = 8'hAE;
        8'd123: galois_lookup_148 = 8'h3A;
        8'd124: galois_lookup_148 = 8'h50;
        8'd125: galois_lookup_148 = 8'hC4;
        8'd126: galois_lookup_148 = 8'hBB;
        8'd127: galois_lookup_148 = 8'h2F;
        8'd128: galois_lookup_148 = 8'hE5;
        8'd129: galois_lookup_148 = 8'h71;
        8'd130: galois_lookup_148 = 8'h0E;
        8'd131: galois_lookup_148 = 8'h9A;
        8'd132: galois_lookup_148 = 8'hF0;
        8'd133: galois_lookup_148 = 8'h64;
        8'd134: galois_lookup_148 = 8'h1B;
        8'd135: galois_lookup_148 = 8'h8F;
        8'd136: galois_lookup_148 = 8'hCF;
        8'd137: galois_lookup_148 = 8'h5B;
        8'd138: galois_lookup_148 = 8'h24;
        8'd139: galois_lookup_148 = 8'hB0;
        8'd140: galois_lookup_148 = 8'hDA;
        8'd141: galois_lookup_148 = 8'h4E;
        8'd142: galois_lookup_148 = 8'h31;
        8'd143: galois_lookup_148 = 8'hA5;
        8'd144: galois_lookup_148 = 8'hB1;
        8'd145: galois_lookup_148 = 8'h25;
        8'd146: galois_lookup_148 = 8'h5A;
        8'd147: galois_lookup_148 = 8'hCE;
        8'd148: galois_lookup_148 = 8'hA4;
        8'd149: galois_lookup_148 = 8'h30;
        8'd150: galois_lookup_148 = 8'h4F;
        8'd151: galois_lookup_148 = 8'hDB;
        8'd152: galois_lookup_148 = 8'h9B;
        8'd153: galois_lookup_148 = 8'h0F;
        8'd154: galois_lookup_148 = 8'h70;
        8'd155: galois_lookup_148 = 8'hE4;
        8'd156: galois_lookup_148 = 8'h8E;
        8'd157: galois_lookup_148 = 8'h1A;
        8'd158: galois_lookup_148 = 8'h65;
        8'd159: galois_lookup_148 = 8'hF1;
        8'd160: galois_lookup_148 = 8'h4D;
        8'd161: galois_lookup_148 = 8'hD9;
        8'd162: galois_lookup_148 = 8'hA6;
        8'd163: galois_lookup_148 = 8'h32;
        8'd164: galois_lookup_148 = 8'h58;
        8'd165: galois_lookup_148 = 8'hCC;
        8'd166: galois_lookup_148 = 8'hB3;
        8'd167: galois_lookup_148 = 8'h27;
        8'd168: galois_lookup_148 = 8'h67;
        8'd169: galois_lookup_148 = 8'hF3;
        8'd170: galois_lookup_148 = 8'h8C;
        8'd171: galois_lookup_148 = 8'h18;
        8'd172: galois_lookup_148 = 8'h72;
        8'd173: galois_lookup_148 = 8'hE6;
        8'd174: galois_lookup_148 = 8'h99;
        8'd175: galois_lookup_148 = 8'h0D;
        8'd176: galois_lookup_148 = 8'h19;
        8'd177: galois_lookup_148 = 8'h8D;
        8'd178: galois_lookup_148 = 8'hF2;
        8'd179: galois_lookup_148 = 8'h66;
        8'd180: galois_lookup_148 = 8'h0C;
        8'd181: galois_lookup_148 = 8'h98;
        8'd182: galois_lookup_148 = 8'hE7;
        8'd183: galois_lookup_148 = 8'h73;
        8'd184: galois_lookup_148 = 8'h33;
        8'd185: galois_lookup_148 = 8'hA7;
        8'd186: galois_lookup_148 = 8'hD8;
        8'd187: galois_lookup_148 = 8'h4C;
        8'd188: galois_lookup_148 = 8'h26;
        8'd189: galois_lookup_148 = 8'hB2;
        8'd190: galois_lookup_148 = 8'hCD;
        8'd191: galois_lookup_148 = 8'h59;
        8'd192: galois_lookup_148 = 8'h76;
        8'd193: galois_lookup_148 = 8'hE2;
        8'd194: galois_lookup_148 = 8'h9D;
        8'd195: galois_lookup_148 = 8'h09;
        8'd196: galois_lookup_148 = 8'h63;
        8'd197: galois_lookup_148 = 8'hF7;
        8'd198: galois_lookup_148 = 8'h88;
        8'd199: galois_lookup_148 = 8'h1C;
        8'd200: galois_lookup_148 = 8'h5C;
        8'd201: galois_lookup_148 = 8'hC8;
        8'd202: galois_lookup_148 = 8'hB7;
        8'd203: galois_lookup_148 = 8'h23;
        8'd204: galois_lookup_148 = 8'h49;
        8'd205: galois_lookup_148 = 8'hDD;
        8'd206: galois_lookup_148 = 8'hA2;
        8'd207: galois_lookup_148 = 8'h36;
        8'd208: galois_lookup_148 = 8'h22;
        8'd209: galois_lookup_148 = 8'hB6;
        8'd210: galois_lookup_148 = 8'hC9;
        8'd211: galois_lookup_148 = 8'h5D;
        8'd212: galois_lookup_148 = 8'h37;
        8'd213: galois_lookup_148 = 8'hA3;
        8'd214: galois_lookup_148 = 8'hDC;
        8'd215: galois_lookup_148 = 8'h48;
        8'd216: galois_lookup_148 = 8'h08;
        8'd217: galois_lookup_148 = 8'h9C;
        8'd218: galois_lookup_148 = 8'hE3;
        8'd219: galois_lookup_148 = 8'h77;
        8'd220: galois_lookup_148 = 8'h1D;
        8'd221: galois_lookup_148 = 8'h89;
        8'd222: galois_lookup_148 = 8'hF6;
        8'd223: galois_lookup_148 = 8'h62;
        8'd224: galois_lookup_148 = 8'hDE;
        8'd225: galois_lookup_148 = 8'h4A;
        8'd226: galois_lookup_148 = 8'h35;
        8'd227: galois_lookup_148 = 8'hA1;
        8'd228: galois_lookup_148 = 8'hCB;
        8'd229: galois_lookup_148 = 8'h5F;
        8'd230: galois_lookup_148 = 8'h20;
        8'd231: galois_lookup_148 = 8'hB4;
        8'd232: galois_lookup_148 = 8'hF4;
        8'd233: galois_lookup_148 = 8'h60;
        8'd234: galois_lookup_148 = 8'h1F;
        8'd235: galois_lookup_148 = 8'h8B;
        8'd236: galois_lookup_148 = 8'hE1;
        8'd237: galois_lookup_148 = 8'h75;
        8'd238: galois_lookup_148 = 8'h0A;
        8'd239: galois_lookup_148 = 8'h9E;
        8'd240: galois_lookup_148 = 8'h8A;
        8'd241: galois_lookup_148 = 8'h1E;
        8'd242: galois_lookup_148 = 8'h61;
        8'd243: galois_lookup_148 = 8'hF5;
        8'd244: galois_lookup_148 = 8'h9F;
        8'd245: galois_lookup_148 = 8'h0B;
        8'd246: galois_lookup_148 = 8'h74;
        8'd247: galois_lookup_148 = 8'hE0;
        8'd248: galois_lookup_148 = 8'hA0;
        8'd249: galois_lookup_148 = 8'h34;
        8'd250: galois_lookup_148 = 8'h4B;
        8'd251: galois_lookup_148 = 8'hDF;
        8'd252: galois_lookup_148 = 8'hB5;
        8'd253: galois_lookup_148 = 8'h21;
        8'd254: galois_lookup_148 = 8'h5E;
        8'd255: galois_lookup_148 = 8'hCA;
    endcase end
endfunction

// -----------------------------------------------------------------------------
function automatic [7:0] galois_lookup_192;
/*

*/
    input   [7:0]   byte;

    begin case (byte)
        8'd000: galois_lookup_192 = 8'h00;
        8'd001: galois_lookup_192 = 8'hC0;
        8'd002: galois_lookup_192 = 8'h43;
        8'd003: galois_lookup_192 = 8'h83;
        8'd004: galois_lookup_192 = 8'h86;
        8'd005: galois_lookup_192 = 8'h46;
        8'd006: galois_lookup_192 = 8'hC5;
        8'd007: galois_lookup_192 = 8'h05;
        8'd008: galois_lookup_192 = 8'hCF;
        8'd009: galois_lookup_192 = 8'h0F;
        8'd010: galois_lookup_192 = 8'h8C;
        8'd011: galois_lookup_192 = 8'h4C;
        8'd012: galois_lookup_192 = 8'h49;
        8'd013: galois_lookup_192 = 8'h89;
        8'd014: galois_lookup_192 = 8'h0A;
        8'd015: galois_lookup_192 = 8'hCA;
        8'd016: galois_lookup_192 = 8'h5D;
        8'd017: galois_lookup_192 = 8'h9D;
        8'd018: galois_lookup_192 = 8'h1E;
        8'd019: galois_lookup_192 = 8'hDE;
        8'd020: galois_lookup_192 = 8'hDB;
        8'd021: galois_lookup_192 = 8'h1B;
        8'd022: galois_lookup_192 = 8'h98;
        8'd023: galois_lookup_192 = 8'h58;
        8'd024: galois_lookup_192 = 8'h92;
        8'd025: galois_lookup_192 = 8'h52;
        8'd026: galois_lookup_192 = 8'hD1;
        8'd027: galois_lookup_192 = 8'h11;
        8'd028: galois_lookup_192 = 8'h14;
        8'd029: galois_lookup_192 = 8'hD4;
        8'd030: galois_lookup_192 = 8'h57;
        8'd031: galois_lookup_192 = 8'h97;
        8'd032: galois_lookup_192 = 8'hBA;
        8'd033: galois_lookup_192 = 8'h7A;
        8'd034: galois_lookup_192 = 8'hF9;
        8'd035: galois_lookup_192 = 8'h39;
        8'd036: galois_lookup_192 = 8'h3C;
        8'd037: galois_lookup_192 = 8'hFC;
        8'd038: galois_lookup_192 = 8'h7F;
        8'd039: galois_lookup_192 = 8'hBF;
        8'd040: galois_lookup_192 = 8'h75;
        8'd041: galois_lookup_192 = 8'hB5;
        8'd042: galois_lookup_192 = 8'h36;
        8'd043: galois_lookup_192 = 8'hF6;
        8'd044: galois_lookup_192 = 8'hF3;
        8'd045: galois_lookup_192 = 8'h33;
        8'd046: galois_lookup_192 = 8'hB0;
        8'd047: galois_lookup_192 = 8'h70;
        8'd048: galois_lookup_192 = 8'hE7;
        8'd049: galois_lookup_192 = 8'h27;
        8'd050: galois_lookup_192 = 8'hA4;
        8'd051: galois_lookup_192 = 8'h64;
        8'd052: galois_lookup_192 = 8'h61;
        8'd053: galois_lookup_192 = 8'hA1;
        8'd054: galois_lookup_192 = 8'h22;
        8'd055: galois_lookup_192 = 8'hE2;
        8'd056: galois_lookup_192 = 8'h28;
        8'd057: galois_lookup_192 = 8'hE8;
        8'd058: galois_lookup_192 = 8'h6B;
        8'd059: galois_lookup_192 = 8'hAB;
        8'd060: galois_lookup_192 = 8'hAE;
        8'd061: galois_lookup_192 = 8'h6E;
        8'd062: galois_lookup_192 = 8'hED;
        8'd063: galois_lookup_192 = 8'h2D;
        8'd064: galois_lookup_192 = 8'hB7;
        8'd065: galois_lookup_192 = 8'h77;
        8'd066: galois_lookup_192 = 8'hF4;
        8'd067: galois_lookup_192 = 8'h34;
        8'd068: galois_lookup_192 = 8'h31;
        8'd069: galois_lookup_192 = 8'hF1;
        8'd070: galois_lookup_192 = 8'h72;
        8'd071: galois_lookup_192 = 8'hB2;
        8'd072: galois_lookup_192 = 8'h78;
        8'd073: galois_lookup_192 = 8'hB8;
        8'd074: galois_lookup_192 = 8'h3B;
        8'd075: galois_lookup_192 = 8'hFB;
        8'd076: galois_lookup_192 = 8'hFE;
        8'd077: galois_lookup_192 = 8'h3E;
        8'd078: galois_lookup_192 = 8'hBD;
        8'd079: galois_lookup_192 = 8'h7D;
        8'd080: galois_lookup_192 = 8'hEA;
        8'd081: galois_lookup_192 = 8'h2A;
        8'd082: galois_lookup_192 = 8'hA9;
        8'd083: galois_lookup_192 = 8'h69;
        8'd084: galois_lookup_192 = 8'h6C;
        8'd085: galois_lookup_192 = 8'hAC;
        8'd086: galois_lookup_192 = 8'h2F;
        8'd087: galois_lookup_192 = 8'hEF;
        8'd088: galois_lookup_192 = 8'h25;
        8'd089: galois_lookup_192 = 8'hE5;
        8'd090: galois_lookup_192 = 8'h66;
        8'd091: galois_lookup_192 = 8'hA6;
        8'd092: galois_lookup_192 = 8'hA3;
        8'd093: galois_lookup_192 = 8'h63;
        8'd094: galois_lookup_192 = 8'hE0;
        8'd095: galois_lookup_192 = 8'h20;
        8'd096: galois_lookup_192 = 8'h0D;
        8'd097: galois_lookup_192 = 8'hCD;
        8'd098: galois_lookup_192 = 8'h4E;
        8'd099: galois_lookup_192 = 8'h8E;
        8'd100: galois_lookup_192 = 8'h8B;
        8'd101: galois_lookup_192 = 8'h4B;
        8'd102: galois_lookup_192 = 8'hC8;
        8'd103: galois_lookup_192 = 8'h08;
        8'd104: galois_lookup_192 = 8'hC2;
        8'd105: galois_lookup_192 = 8'h02;
        8'd106: galois_lookup_192 = 8'h81;
        8'd107: galois_lookup_192 = 8'h41;
        8'd108: galois_lookup_192 = 8'h44;
        8'd109: galois_lookup_192 = 8'h84;
        8'd110: galois_lookup_192 = 8'h07;
        8'd111: galois_lookup_192 = 8'hC7;
        8'd112: galois_lookup_192 = 8'h50;
        8'd113: galois_lookup_192 = 8'h90;
        8'd114: galois_lookup_192 = 8'h13;
        8'd115: galois_lookup_192 = 8'hD3;
        8'd116: galois_lookup_192 = 8'hD6;
        8'd117: galois_lookup_192 = 8'h16;
        8'd118: galois_lookup_192 = 8'h95;
        8'd119: galois_lookup_192 = 8'h55;
        8'd120: galois_lookup_192 = 8'h9F;
        8'd121: galois_lookup_192 = 8'h5F;
        8'd122: galois_lookup_192 = 8'hDC;
        8'd123: galois_lookup_192 = 8'h1C;
        8'd124: galois_lookup_192 = 8'h19;
        8'd125: galois_lookup_192 = 8'hD9;
        8'd126: galois_lookup_192 = 8'h5A;
        8'd127: galois_lookup_192 = 8'h9A;
        8'd128: galois_lookup_192 = 8'hAD;
        8'd129: galois_lookup_192 = 8'h6D;
        8'd130: galois_lookup_192 = 8'hEE;
        8'd131: galois_lookup_192 = 8'h2E;
        8'd132: galois_lookup_192 = 8'h2B;
        8'd133: galois_lookup_192 = 8'hEB;
        8'd134: galois_lookup_192 = 8'h68;
        8'd135: galois_lookup_192 = 8'hA8;
        8'd136: galois_lookup_192 = 8'h62;
        8'd137: galois_lookup_192 = 8'hA2;
        8'd138: galois_lookup_192 = 8'h21;
        8'd139: galois_lookup_192 = 8'hE1;
        8'd140: galois_lookup_192 = 8'hE4;
        8'd141: galois_lookup_192 = 8'h24;
        8'd142: galois_lookup_192 = 8'hA7;
        8'd143: galois_lookup_192 = 8'h67;
        8'd144: galois_lookup_192 = 8'hF0;
        8'd145: galois_lookup_192 = 8'h30;
        8'd146: galois_lookup_192 = 8'hB3;
        8'd147: galois_lookup_192 = 8'h73;
        8'd148: galois_lookup_192 = 8'h76;
        8'd149: galois_lookup_192 = 8'hB6;
        8'd150: galois_lookup_192 = 8'h35;
        8'd151: galois_lookup_192 = 8'hF5;
        8'd152: galois_lookup_192 = 8'h3F;
        8'd153: galois_lookup_192 = 8'hFF;
        8'd154: galois_lookup_192 = 8'h7C;
        8'd155: galois_lookup_192 = 8'hBC;
        8'd156: galois_lookup_192 = 8'hB9;
        8'd157: galois_lookup_192 = 8'h79;
        8'd158: galois_lookup_192 = 8'hFA;
        8'd159: galois_lookup_192 = 8'h3A;
        8'd160: galois_lookup_192 = 8'h17;
        8'd161: galois_lookup_192 = 8'hD7;
        8'd162: galois_lookup_192 = 8'h54;
        8'd163: galois_lookup_192 = 8'h94;
        8'd164: galois_lookup_192 = 8'h91;
        8'd165: galois_lookup_192 = 8'h51;
        8'd166: galois_lookup_192 = 8'hD2;
        8'd167: galois_lookup_192 = 8'h12;
        8'd168: galois_lookup_192 = 8'hD8;
        8'd169: galois_lookup_192 = 8'h18;
        8'd170: galois_lookup_192 = 8'h9B;
        8'd171: galois_lookup_192 = 8'h5B;
        8'd172: galois_lookup_192 = 8'h5E;
        8'd173: galois_lookup_192 = 8'h9E;
        8'd174: galois_lookup_192 = 8'h1D;
        8'd175: galois_lookup_192 = 8'hDD;
        8'd176: galois_lookup_192 = 8'h4A;
        8'd177: galois_lookup_192 = 8'h8A;
        8'd178: galois_lookup_192 = 8'h09;
        8'd179: galois_lookup_192 = 8'hC9;
        8'd180: galois_lookup_192 = 8'hCC;
        8'd181: galois_lookup_192 = 8'h0C;
        8'd182: galois_lookup_192 = 8'h8F;
        8'd183: galois_lookup_192 = 8'h4F;
        8'd184: galois_lookup_192 = 8'h85;
        8'd185: galois_lookup_192 = 8'h45;
        8'd186: galois_lookup_192 = 8'hC6;
        8'd187: galois_lookup_192 = 8'h06;
        8'd188: galois_lookup_192 = 8'h03;
        8'd189: galois_lookup_192 = 8'hC3;
        8'd190: galois_lookup_192 = 8'h40;
        8'd191: galois_lookup_192 = 8'h80;
        8'd192: galois_lookup_192 = 8'h1A;
        8'd193: galois_lookup_192 = 8'hDA;
        8'd194: galois_lookup_192 = 8'h59;
        8'd195: galois_lookup_192 = 8'h99;
        8'd196: galois_lookup_192 = 8'h9C;
        8'd197: galois_lookup_192 = 8'h5C;
        8'd198: galois_lookup_192 = 8'hDF;
        8'd199: galois_lookup_192 = 8'h1F;
        8'd200: galois_lookup_192 = 8'hD5;
        8'd201: galois_lookup_192 = 8'h15;
        8'd202: galois_lookup_192 = 8'h96;
        8'd203: galois_lookup_192 = 8'h56;
        8'd204: galois_lookup_192 = 8'h53;
        8'd205: galois_lookup_192 = 8'h93;
        8'd206: galois_lookup_192 = 8'h10;
        8'd207: galois_lookup_192 = 8'hD0;
        8'd208: galois_lookup_192 = 8'h47;
        8'd209: galois_lookup_192 = 8'h87;
        8'd210: galois_lookup_192 = 8'h04;
        8'd211: galois_lookup_192 = 8'hC4;
        8'd212: galois_lookup_192 = 8'hC1;
        8'd213: galois_lookup_192 = 8'h01;
        8'd214: galois_lookup_192 = 8'h82;
        8'd215: galois_lookup_192 = 8'h42;
        8'd216: galois_lookup_192 = 8'h88;
        8'd217: galois_lookup_192 = 8'h48;
        8'd218: galois_lookup_192 = 8'hCB;
        8'd219: galois_lookup_192 = 8'h0B;
        8'd220: galois_lookup_192 = 8'h0E;
        8'd221: galois_lookup_192 = 8'hCE;
        8'd222: galois_lookup_192 = 8'h4D;
        8'd223: galois_lookup_192 = 8'h8D;
        8'd224: galois_lookup_192 = 8'hA0;
        8'd225: galois_lookup_192 = 8'h60;
        8'd226: galois_lookup_192 = 8'hE3;
        8'd227: galois_lookup_192 = 8'h23;
        8'd228: galois_lookup_192 = 8'h26;
        8'd229: galois_lookup_192 = 8'hE6;
        8'd230: galois_lookup_192 = 8'h65;
        8'd231: galois_lookup_192 = 8'hA5;
        8'd232: galois_lookup_192 = 8'h6F;
        8'd233: galois_lookup_192 = 8'hAF;
        8'd234: galois_lookup_192 = 8'h2C;
        8'd235: galois_lookup_192 = 8'hEC;
        8'd236: galois_lookup_192 = 8'hE9;
        8'd237: galois_lookup_192 = 8'h29;
        8'd238: galois_lookup_192 = 8'hAA;
        8'd239: galois_lookup_192 = 8'h6A;
        8'd240: galois_lookup_192 = 8'hFD;
        8'd241: galois_lookup_192 = 8'h3D;
        8'd242: galois_lookup_192 = 8'hBE;
        8'd243: galois_lookup_192 = 8'h7E;
        8'd244: galois_lookup_192 = 8'h7B;
        8'd245: galois_lookup_192 = 8'hBB;
        8'd246: galois_lookup_192 = 8'h38;
        8'd247: galois_lookup_192 = 8'hF8;
        8'd248: galois_lookup_192 = 8'h32;
        8'd249: galois_lookup_192 = 8'hF2;
        8'd250: galois_lookup_192 = 8'h71;
        8'd251: galois_lookup_192 = 8'hB1;
        8'd252: galois_lookup_192 = 8'hB4;
        8'd253: galois_lookup_192 = 8'h74;
        8'd254: galois_lookup_192 = 8'hF7;
        8'd255: galois_lookup_192 = 8'h37;
    endcase end
endfunction

// -----------------------------------------------------------------------------
function automatic [7:0] galois_lookup_194;
/*

*/
    input   [7:0]   byte;

    begin case (byte)
        8'd000: galois_lookup_194 = 8'h00;
        8'd001: galois_lookup_194 = 8'hC2;
        8'd002: galois_lookup_194 = 8'h47;
        8'd003: galois_lookup_194 = 8'h85;
        8'd004: galois_lookup_194 = 8'h8E;
        8'd005: galois_lookup_194 = 8'h4C;
        8'd006: galois_lookup_194 = 8'hC9;
        8'd007: galois_lookup_194 = 8'h0B;
        8'd008: galois_lookup_194 = 8'hDF;
        8'd009: galois_lookup_194 = 8'h1D;
        8'd010: galois_lookup_194 = 8'h98;
        8'd011: galois_lookup_194 = 8'h5A;
        8'd012: galois_lookup_194 = 8'h51;
        8'd013: galois_lookup_194 = 8'h93;
        8'd014: galois_lookup_194 = 8'h16;
        8'd015: galois_lookup_194 = 8'hD4;
        8'd016: galois_lookup_194 = 8'h7D;
        8'd017: galois_lookup_194 = 8'hBF;
        8'd018: galois_lookup_194 = 8'h3A;
        8'd019: galois_lookup_194 = 8'hF8;
        8'd020: galois_lookup_194 = 8'hF3;
        8'd021: galois_lookup_194 = 8'h31;
        8'd022: galois_lookup_194 = 8'hB4;
        8'd023: galois_lookup_194 = 8'h76;
        8'd024: galois_lookup_194 = 8'hA2;
        8'd025: galois_lookup_194 = 8'h60;
        8'd026: galois_lookup_194 = 8'hE5;
        8'd027: galois_lookup_194 = 8'h27;
        8'd028: galois_lookup_194 = 8'h2C;
        8'd029: galois_lookup_194 = 8'hEE;
        8'd030: galois_lookup_194 = 8'h6B;
        8'd031: galois_lookup_194 = 8'hA9;
        8'd032: galois_lookup_194 = 8'hFA;
        8'd033: galois_lookup_194 = 8'h38;
        8'd034: galois_lookup_194 = 8'hBD;
        8'd035: galois_lookup_194 = 8'h7F;
        8'd036: galois_lookup_194 = 8'h74;
        8'd037: galois_lookup_194 = 8'hB6;
        8'd038: galois_lookup_194 = 8'h33;
        8'd039: galois_lookup_194 = 8'hF1;
        8'd040: galois_lookup_194 = 8'h25;
        8'd041: galois_lookup_194 = 8'hE7;
        8'd042: galois_lookup_194 = 8'h62;
        8'd043: galois_lookup_194 = 8'hA0;
        8'd044: galois_lookup_194 = 8'hAB;
        8'd045: galois_lookup_194 = 8'h69;
        8'd046: galois_lookup_194 = 8'hEC;
        8'd047: galois_lookup_194 = 8'h2E;
        8'd048: galois_lookup_194 = 8'h87;
        8'd049: galois_lookup_194 = 8'h45;
        8'd050: galois_lookup_194 = 8'hC0;
        8'd051: galois_lookup_194 = 8'h02;
        8'd052: galois_lookup_194 = 8'h09;
        8'd053: galois_lookup_194 = 8'hCB;
        8'd054: galois_lookup_194 = 8'h4E;
        8'd055: galois_lookup_194 = 8'h8C;
        8'd056: galois_lookup_194 = 8'h58;
        8'd057: galois_lookup_194 = 8'h9A;
        8'd058: galois_lookup_194 = 8'h1F;
        8'd059: galois_lookup_194 = 8'hDD;
        8'd060: galois_lookup_194 = 8'hD6;
        8'd061: galois_lookup_194 = 8'h14;
        8'd062: galois_lookup_194 = 8'h91;
        8'd063: galois_lookup_194 = 8'h53;
        8'd064: galois_lookup_194 = 8'h37;
        8'd065: galois_lookup_194 = 8'hF5;
        8'd066: galois_lookup_194 = 8'h70;
        8'd067: galois_lookup_194 = 8'hB2;
        8'd068: galois_lookup_194 = 8'hB9;
        8'd069: galois_lookup_194 = 8'h7B;
        8'd070: galois_lookup_194 = 8'hFE;
        8'd071: galois_lookup_194 = 8'h3C;
        8'd072: galois_lookup_194 = 8'hE8;
        8'd073: galois_lookup_194 = 8'h2A;
        8'd074: galois_lookup_194 = 8'hAF;
        8'd075: galois_lookup_194 = 8'h6D;
        8'd076: galois_lookup_194 = 8'h66;
        8'd077: galois_lookup_194 = 8'hA4;
        8'd078: galois_lookup_194 = 8'h21;
        8'd079: galois_lookup_194 = 8'hE3;
        8'd080: galois_lookup_194 = 8'h4A;
        8'd081: galois_lookup_194 = 8'h88;
        8'd082: galois_lookup_194 = 8'h0D;
        8'd083: galois_lookup_194 = 8'hCF;
        8'd084: galois_lookup_194 = 8'hC4;
        8'd085: galois_lookup_194 = 8'h06;
        8'd086: galois_lookup_194 = 8'h83;
        8'd087: galois_lookup_194 = 8'h41;
        8'd088: galois_lookup_194 = 8'h95;
        8'd089: galois_lookup_194 = 8'h57;
        8'd090: galois_lookup_194 = 8'hD2;
        8'd091: galois_lookup_194 = 8'h10;
        8'd092: galois_lookup_194 = 8'h1B;
        8'd093: galois_lookup_194 = 8'hD9;
        8'd094: galois_lookup_194 = 8'h5C;
        8'd095: galois_lookup_194 = 8'h9E;
        8'd096: galois_lookup_194 = 8'hCD;
        8'd097: galois_lookup_194 = 8'h0F;
        8'd098: galois_lookup_194 = 8'h8A;
        8'd099: galois_lookup_194 = 8'h48;
        8'd100: galois_lookup_194 = 8'h43;
        8'd101: galois_lookup_194 = 8'h81;
        8'd102: galois_lookup_194 = 8'h04;
        8'd103: galois_lookup_194 = 8'hC6;
        8'd104: galois_lookup_194 = 8'h12;
        8'd105: galois_lookup_194 = 8'hD0;
        8'd106: galois_lookup_194 = 8'h55;
        8'd107: galois_lookup_194 = 8'h97;
        8'd108: galois_lookup_194 = 8'h9C;
        8'd109: galois_lookup_194 = 8'h5E;
        8'd110: galois_lookup_194 = 8'hDB;
        8'd111: galois_lookup_194 = 8'h19;
        8'd112: galois_lookup_194 = 8'hB0;
        8'd113: galois_lookup_194 = 8'h72;
        8'd114: galois_lookup_194 = 8'hF7;
        8'd115: galois_lookup_194 = 8'h35;
        8'd116: galois_lookup_194 = 8'h3E;
        8'd117: galois_lookup_194 = 8'hFC;
        8'd118: galois_lookup_194 = 8'h79;
        8'd119: galois_lookup_194 = 8'hBB;
        8'd120: galois_lookup_194 = 8'h6F;
        8'd121: galois_lookup_194 = 8'hAD;
        8'd122: galois_lookup_194 = 8'h28;
        8'd123: galois_lookup_194 = 8'hEA;
        8'd124: galois_lookup_194 = 8'hE1;
        8'd125: galois_lookup_194 = 8'h23;
        8'd126: galois_lookup_194 = 8'hA6;
        8'd127: galois_lookup_194 = 8'h64;
        8'd128: galois_lookup_194 = 8'h6E;
        8'd129: galois_lookup_194 = 8'hAC;
        8'd130: galois_lookup_194 = 8'h29;
        8'd131: galois_lookup_194 = 8'hEB;
        8'd132: galois_lookup_194 = 8'hE0;
        8'd133: galois_lookup_194 = 8'h22;
        8'd134: galois_lookup_194 = 8'hA7;
        8'd135: galois_lookup_194 = 8'h65;
        8'd136: galois_lookup_194 = 8'hB1;
        8'd137: galois_lookup_194 = 8'h73;
        8'd138: galois_lookup_194 = 8'hF6;
        8'd139: galois_lookup_194 = 8'h34;
        8'd140: galois_lookup_194 = 8'h3F;
        8'd141: galois_lookup_194 = 8'hFD;
        8'd142: galois_lookup_194 = 8'h78;
        8'd143: galois_lookup_194 = 8'hBA;
        8'd144: galois_lookup_194 = 8'h13;
        8'd145: galois_lookup_194 = 8'hD1;
        8'd146: galois_lookup_194 = 8'h54;
        8'd147: galois_lookup_194 = 8'h96;
        8'd148: galois_lookup_194 = 8'h9D;
        8'd149: galois_lookup_194 = 8'h5F;
        8'd150: galois_lookup_194 = 8'hDA;
        8'd151: galois_lookup_194 = 8'h18;
        8'd152: galois_lookup_194 = 8'hCC;
        8'd153: galois_lookup_194 = 8'h0E;
        8'd154: galois_lookup_194 = 8'h8B;
        8'd155: galois_lookup_194 = 8'h49;
        8'd156: galois_lookup_194 = 8'h42;
        8'd157: galois_lookup_194 = 8'h80;
        8'd158: galois_lookup_194 = 8'h05;
        8'd159: galois_lookup_194 = 8'hC7;
        8'd160: galois_lookup_194 = 8'h94;
        8'd161: galois_lookup_194 = 8'h56;
        8'd162: galois_lookup_194 = 8'hD3;
        8'd163: galois_lookup_194 = 8'h11;
        8'd164: galois_lookup_194 = 8'h1A;
        8'd165: galois_lookup_194 = 8'hD8;
        8'd166: galois_lookup_194 = 8'h5D;
        8'd167: galois_lookup_194 = 8'h9F;
        8'd168: galois_lookup_194 = 8'h4B;
        8'd169: galois_lookup_194 = 8'h89;
        8'd170: galois_lookup_194 = 8'h0C;
        8'd171: galois_lookup_194 = 8'hCE;
        8'd172: galois_lookup_194 = 8'hC5;
        8'd173: galois_lookup_194 = 8'h07;
        8'd174: galois_lookup_194 = 8'h82;
        8'd175: galois_lookup_194 = 8'h40;
        8'd176: galois_lookup_194 = 8'hE9;
        8'd177: galois_lookup_194 = 8'h2B;
        8'd178: galois_lookup_194 = 8'hAE;
        8'd179: galois_lookup_194 = 8'h6C;
        8'd180: galois_lookup_194 = 8'h67;
        8'd181: galois_lookup_194 = 8'hA5;
        8'd182: galois_lookup_194 = 8'h20;
        8'd183: galois_lookup_194 = 8'hE2;
        8'd184: galois_lookup_194 = 8'h36;
        8'd185: galois_lookup_194 = 8'hF4;
        8'd186: galois_lookup_194 = 8'h71;
        8'd187: galois_lookup_194 = 8'hB3;
        8'd188: galois_lookup_194 = 8'hB8;
        8'd189: galois_lookup_194 = 8'h7A;
        8'd190: galois_lookup_194 = 8'hFF;
        8'd191: galois_lookup_194 = 8'h3D;
        8'd192: galois_lookup_194 = 8'h59;
        8'd193: galois_lookup_194 = 8'h9B;
        8'd194: galois_lookup_194 = 8'h1E;
        8'd195: galois_lookup_194 = 8'hDC;
        8'd196: galois_lookup_194 = 8'hD7;
        8'd197: galois_lookup_194 = 8'h15;
        8'd198: galois_lookup_194 = 8'h90;
        8'd199: galois_lookup_194 = 8'h52;
        8'd200: galois_lookup_194 = 8'h86;
        8'd201: galois_lookup_194 = 8'h44;
        8'd202: galois_lookup_194 = 8'hC1;
        8'd203: galois_lookup_194 = 8'h03;
        8'd204: galois_lookup_194 = 8'h08;
        8'd205: galois_lookup_194 = 8'hCA;
        8'd206: galois_lookup_194 = 8'h4F;
        8'd207: galois_lookup_194 = 8'h8D;
        8'd208: galois_lookup_194 = 8'h24;
        8'd209: galois_lookup_194 = 8'hE6;
        8'd210: galois_lookup_194 = 8'h63;
        8'd211: galois_lookup_194 = 8'hA1;
        8'd212: galois_lookup_194 = 8'hAA;
        8'd213: galois_lookup_194 = 8'h68;
        8'd214: galois_lookup_194 = 8'hED;
        8'd215: galois_lookup_194 = 8'h2F;
        8'd216: galois_lookup_194 = 8'hFB;
        8'd217: galois_lookup_194 = 8'h39;
        8'd218: galois_lookup_194 = 8'hBC;
        8'd219: galois_lookup_194 = 8'h7E;
        8'd220: galois_lookup_194 = 8'h75;
        8'd221: galois_lookup_194 = 8'hB7;
        8'd222: galois_lookup_194 = 8'h32;
        8'd223: galois_lookup_194 = 8'hF0;
        8'd224: galois_lookup_194 = 8'hA3;
        8'd225: galois_lookup_194 = 8'h61;
        8'd226: galois_lookup_194 = 8'hE4;
        8'd227: galois_lookup_194 = 8'h26;
        8'd228: galois_lookup_194 = 8'h2D;
        8'd229: galois_lookup_194 = 8'hEF;
        8'd230: galois_lookup_194 = 8'h6A;
        8'd231: galois_lookup_194 = 8'hA8;
        8'd232: galois_lookup_194 = 8'h7C;
        8'd233: galois_lookup_194 = 8'hBE;
        8'd234: galois_lookup_194 = 8'h3B;
        8'd235: galois_lookup_194 = 8'hF9;
        8'd236: galois_lookup_194 = 8'hF2;
        8'd237: galois_lookup_194 = 8'h30;
        8'd238: galois_lookup_194 = 8'hB5;
        8'd239: galois_lookup_194 = 8'h77;
        8'd240: galois_lookup_194 = 8'hDE;
        8'd241: galois_lookup_194 = 8'h1C;
        8'd242: galois_lookup_194 = 8'h99;
        8'd243: galois_lookup_194 = 8'h5B;
        8'd244: galois_lookup_194 = 8'h50;
        8'd245: galois_lookup_194 = 8'h92;
        8'd246: galois_lookup_194 = 8'h17;
        8'd247: galois_lookup_194 = 8'hD5;
        8'd248: galois_lookup_194 = 8'h01;
        8'd249: galois_lookup_194 = 8'hC3;
        8'd250: galois_lookup_194 = 8'h46;
        8'd251: galois_lookup_194 = 8'h84;
        8'd252: galois_lookup_194 = 8'h8F;
        8'd253: galois_lookup_194 = 8'h4D;
        8'd254: galois_lookup_194 = 8'hC8;
        8'd255: galois_lookup_194 = 8'h0A;
    endcase end
endfunction

// -----------------------------------------------------------------------------
function automatic [7:0] galois_lookup_251;
/*

*/
    input   [7:0]   byte;

    begin case (byte)
        8'd000: galois_lookup_251 = 8'h00;
        8'd001: galois_lookup_251 = 8'hFB;
        8'd002: galois_lookup_251 = 8'h35;
        8'd003: galois_lookup_251 = 8'hCE;
        8'd004: galois_lookup_251 = 8'h6A;
        8'd005: galois_lookup_251 = 8'h91;
        8'd006: galois_lookup_251 = 8'h5F;
        8'd007: galois_lookup_251 = 8'hA4;
        8'd008: galois_lookup_251 = 8'hD4;
        8'd009: galois_lookup_251 = 8'h2F;
        8'd010: galois_lookup_251 = 8'hE1;
        8'd011: galois_lookup_251 = 8'h1A;
        8'd012: galois_lookup_251 = 8'hBE;
        8'd013: galois_lookup_251 = 8'h45;
        8'd014: galois_lookup_251 = 8'h8B;
        8'd015: galois_lookup_251 = 8'h70;
        8'd016: galois_lookup_251 = 8'h6B;
        8'd017: galois_lookup_251 = 8'h90;
        8'd018: galois_lookup_251 = 8'h5E;
        8'd019: galois_lookup_251 = 8'hA5;
        8'd020: galois_lookup_251 = 8'h01;
        8'd021: galois_lookup_251 = 8'hFA;
        8'd022: galois_lookup_251 = 8'h34;
        8'd023: galois_lookup_251 = 8'hCF;
        8'd024: galois_lookup_251 = 8'hBF;
        8'd025: galois_lookup_251 = 8'h44;
        8'd026: galois_lookup_251 = 8'h8A;
        8'd027: galois_lookup_251 = 8'h71;
        8'd028: galois_lookup_251 = 8'hD5;
        8'd029: galois_lookup_251 = 8'h2E;
        8'd030: galois_lookup_251 = 8'hE0;
        8'd031: galois_lookup_251 = 8'h1B;
        8'd032: galois_lookup_251 = 8'hD6;
        8'd033: galois_lookup_251 = 8'h2D;
        8'd034: galois_lookup_251 = 8'hE3;
        8'd035: galois_lookup_251 = 8'h18;
        8'd036: galois_lookup_251 = 8'hBC;
        8'd037: galois_lookup_251 = 8'h47;
        8'd038: galois_lookup_251 = 8'h89;
        8'd039: galois_lookup_251 = 8'h72;
        8'd040: galois_lookup_251 = 8'h02;
        8'd041: galois_lookup_251 = 8'hF9;
        8'd042: galois_lookup_251 = 8'h37;
        8'd043: galois_lookup_251 = 8'hCC;
        8'd044: galois_lookup_251 = 8'h68;
        8'd045: galois_lookup_251 = 8'h93;
        8'd046: galois_lookup_251 = 8'h5D;
        8'd047: galois_lookup_251 = 8'hA6;
        8'd048: galois_lookup_251 = 8'hBD;
        8'd049: galois_lookup_251 = 8'h46;
        8'd050: galois_lookup_251 = 8'h88;
        8'd051: galois_lookup_251 = 8'h73;
        8'd052: galois_lookup_251 = 8'hD7;
        8'd053: galois_lookup_251 = 8'h2C;
        8'd054: galois_lookup_251 = 8'hE2;
        8'd055: galois_lookup_251 = 8'h19;
        8'd056: galois_lookup_251 = 8'h69;
        8'd057: galois_lookup_251 = 8'h92;
        8'd058: galois_lookup_251 = 8'h5C;
        8'd059: galois_lookup_251 = 8'hA7;
        8'd060: galois_lookup_251 = 8'h03;
        8'd061: galois_lookup_251 = 8'hF8;
        8'd062: galois_lookup_251 = 8'h36;
        8'd063: galois_lookup_251 = 8'hCD;
        8'd064: galois_lookup_251 = 8'h6F;
        8'd065: galois_lookup_251 = 8'h94;
        8'd066: galois_lookup_251 = 8'h5A;
        8'd067: galois_lookup_251 = 8'hA1;
        8'd068: galois_lookup_251 = 8'h05;
        8'd069: galois_lookup_251 = 8'hFE;
        8'd070: galois_lookup_251 = 8'h30;
        8'd071: galois_lookup_251 = 8'hCB;
        8'd072: galois_lookup_251 = 8'hBB;
        8'd073: galois_lookup_251 = 8'h40;
        8'd074: galois_lookup_251 = 8'h8E;
        8'd075: galois_lookup_251 = 8'h75;
        8'd076: galois_lookup_251 = 8'hD1;
        8'd077: galois_lookup_251 = 8'h2A;
        8'd078: galois_lookup_251 = 8'hE4;
        8'd079: galois_lookup_251 = 8'h1F;
        8'd080: galois_lookup_251 = 8'h04;
        8'd081: galois_lookup_251 = 8'hFF;
        8'd082: galois_lookup_251 = 8'h31;
        8'd083: galois_lookup_251 = 8'hCA;
        8'd084: galois_lookup_251 = 8'h6E;
        8'd085: galois_lookup_251 = 8'h95;
        8'd086: galois_lookup_251 = 8'h5B;
        8'd087: galois_lookup_251 = 8'hA0;
        8'd088: galois_lookup_251 = 8'hD0;
        8'd089: galois_lookup_251 = 8'h2B;
        8'd090: galois_lookup_251 = 8'hE5;
        8'd091: galois_lookup_251 = 8'h1E;
        8'd092: galois_lookup_251 = 8'hBA;
        8'd093: galois_lookup_251 = 8'h41;
        8'd094: galois_lookup_251 = 8'h8F;
        8'd095: galois_lookup_251 = 8'h74;
        8'd096: galois_lookup_251 = 8'hB9;
        8'd097: galois_lookup_251 = 8'h42;
        8'd098: galois_lookup_251 = 8'h8C;
        8'd099: galois_lookup_251 = 8'h77;
        8'd100: galois_lookup_251 = 8'hD3;
        8'd101: galois_lookup_251 = 8'h28;
        8'd102: galois_lookup_251 = 8'hE6;
        8'd103: galois_lookup_251 = 8'h1D;
        8'd104: galois_lookup_251 = 8'h6D;
        8'd105: galois_lookup_251 = 8'h96;
        8'd106: galois_lookup_251 = 8'h58;
        8'd107: galois_lookup_251 = 8'hA3;
        8'd108: galois_lookup_251 = 8'h07;
        8'd109: galois_lookup_251 = 8'hFC;
        8'd110: galois_lookup_251 = 8'h32;
        8'd111: galois_lookup_251 = 8'hC9;
        8'd112: galois_lookup_251 = 8'hD2;
        8'd113: galois_lookup_251 = 8'h29;
        8'd114: galois_lookup_251 = 8'hE7;
        8'd115: galois_lookup_251 = 8'h1C;
        8'd116: galois_lookup_251 = 8'hB8;
        8'd117: galois_lookup_251 = 8'h43;
        8'd118: galois_lookup_251 = 8'h8D;
        8'd119: galois_lookup_251 = 8'h76;
        8'd120: galois_lookup_251 = 8'h06;
        8'd121: galois_lookup_251 = 8'hFD;
        8'd122: galois_lookup_251 = 8'h33;
        8'd123: galois_lookup_251 = 8'hC8;
        8'd124: galois_lookup_251 = 8'h6C;
        8'd125: galois_lookup_251 = 8'h97;
        8'd126: galois_lookup_251 = 8'h59;
        8'd127: galois_lookup_251 = 8'hA2;
        8'd128: galois_lookup_251 = 8'hDE;
        8'd129: galois_lookup_251 = 8'h25;
        8'd130: galois_lookup_251 = 8'hEB;
        8'd131: galois_lookup_251 = 8'h10;
        8'd132: galois_lookup_251 = 8'hB4;
        8'd133: galois_lookup_251 = 8'h4F;
        8'd134: galois_lookup_251 = 8'h81;
        8'd135: galois_lookup_251 = 8'h7A;
        8'd136: galois_lookup_251 = 8'h0A;
        8'd137: galois_lookup_251 = 8'hF1;
        8'd138: galois_lookup_251 = 8'h3F;
        8'd139: galois_lookup_251 = 8'hC4;
        8'd140: galois_lookup_251 = 8'h60;
        8'd141: galois_lookup_251 = 8'h9B;
        8'd142: galois_lookup_251 = 8'h55;
        8'd143: galois_lookup_251 = 8'hAE;
        8'd144: galois_lookup_251 = 8'hB5;
        8'd145: galois_lookup_251 = 8'h4E;
        8'd146: galois_lookup_251 = 8'h80;
        8'd147: galois_lookup_251 = 8'h7B;
        8'd148: galois_lookup_251 = 8'hDF;
        8'd149: galois_lookup_251 = 8'h24;
        8'd150: galois_lookup_251 = 8'hEA;
        8'd151: galois_lookup_251 = 8'h11;
        8'd152: galois_lookup_251 = 8'h61;
        8'd153: galois_lookup_251 = 8'h9A;
        8'd154: galois_lookup_251 = 8'h54;
        8'd155: galois_lookup_251 = 8'hAF;
        8'd156: galois_lookup_251 = 8'h0B;
        8'd157: galois_lookup_251 = 8'hF0;
        8'd158: galois_lookup_251 = 8'h3E;
        8'd159: galois_lookup_251 = 8'hC5;
        8'd160: galois_lookup_251 = 8'h08;
        8'd161: galois_lookup_251 = 8'hF3;
        8'd162: galois_lookup_251 = 8'h3D;
        8'd163: galois_lookup_251 = 8'hC6;
        8'd164: galois_lookup_251 = 8'h62;
        8'd165: galois_lookup_251 = 8'h99;
        8'd166: galois_lookup_251 = 8'h57;
        8'd167: galois_lookup_251 = 8'hAC;
        8'd168: galois_lookup_251 = 8'hDC;
        8'd169: galois_lookup_251 = 8'h27;
        8'd170: galois_lookup_251 = 8'hE9;
        8'd171: galois_lookup_251 = 8'h12;
        8'd172: galois_lookup_251 = 8'hB6;
        8'd173: galois_lookup_251 = 8'h4D;
        8'd174: galois_lookup_251 = 8'h83;
        8'd175: galois_lookup_251 = 8'h78;
        8'd176: galois_lookup_251 = 8'h63;
        8'd177: galois_lookup_251 = 8'h98;
        8'd178: galois_lookup_251 = 8'h56;
        8'd179: galois_lookup_251 = 8'hAD;
        8'd180: galois_lookup_251 = 8'h09;
        8'd181: galois_lookup_251 = 8'hF2;
        8'd182: galois_lookup_251 = 8'h3C;
        8'd183: galois_lookup_251 = 8'hC7;
        8'd184: galois_lookup_251 = 8'hB7;
        8'd185: galois_lookup_251 = 8'h4C;
        8'd186: galois_lookup_251 = 8'h82;
        8'd187: galois_lookup_251 = 8'h79;
        8'd188: galois_lookup_251 = 8'hDD;
        8'd189: galois_lookup_251 = 8'h26;
        8'd190: galois_lookup_251 = 8'hE8;
        8'd191: galois_lookup_251 = 8'h13;
        8'd192: galois_lookup_251 = 8'hB1;
        8'd193: galois_lookup_251 = 8'h4A;
        8'd194: galois_lookup_251 = 8'h84;
        8'd195: galois_lookup_251 = 8'h7F;
        8'd196: galois_lookup_251 = 8'hDB;
        8'd197: galois_lookup_251 = 8'h20;
        8'd198: galois_lookup_251 = 8'hEE;
        8'd199: galois_lookup_251 = 8'h15;
        8'd200: galois_lookup_251 = 8'h65;
        8'd201: galois_lookup_251 = 8'h9E;
        8'd202: galois_lookup_251 = 8'h50;
        8'd203: galois_lookup_251 = 8'hAB;
        8'd204: galois_lookup_251 = 8'h0F;
        8'd205: galois_lookup_251 = 8'hF4;
        8'd206: galois_lookup_251 = 8'h3A;
        8'd207: galois_lookup_251 = 8'hC1;
        8'd208: galois_lookup_251 = 8'hDA;
        8'd209: galois_lookup_251 = 8'h21;
        8'd210: galois_lookup_251 = 8'hEF;
        8'd211: galois_lookup_251 = 8'h14;
        8'd212: galois_lookup_251 = 8'hB0;
        8'd213: galois_lookup_251 = 8'h4B;
        8'd214: galois_lookup_251 = 8'h85;
        8'd215: galois_lookup_251 = 8'h7E;
        8'd216: galois_lookup_251 = 8'h0E;
        8'd217: galois_lookup_251 = 8'hF5;
        8'd218: galois_lookup_251 = 8'h3B;
        8'd219: galois_lookup_251 = 8'hC0;
        8'd220: galois_lookup_251 = 8'h64;
        8'd221: galois_lookup_251 = 8'h9F;
        8'd222: galois_lookup_251 = 8'h51;
        8'd223: galois_lookup_251 = 8'hAA;
        8'd224: galois_lookup_251 = 8'h67;
        8'd225: galois_lookup_251 = 8'h9C;
        8'd226: galois_lookup_251 = 8'h52;
        8'd227: galois_lookup_251 = 8'hA9;
        8'd228: galois_lookup_251 = 8'h0D;
        8'd229: galois_lookup_251 = 8'hF6;
        8'd230: galois_lookup_251 = 8'h38;
        8'd231: galois_lookup_251 = 8'hC3;
        8'd232: galois_lookup_251 = 8'hB3;
        8'd233: galois_lookup_251 = 8'h48;
        8'd234: galois_lookup_251 = 8'h86;
        8'd235: galois_lookup_251 = 8'h7D;
        8'd236: galois_lookup_251 = 8'hD9;
        8'd237: galois_lookup_251 = 8'h22;
        8'd238: galois_lookup_251 = 8'hEC;
        8'd239: galois_lookup_251 = 8'h17;
        8'd240: galois_lookup_251 = 8'h0C;
        8'd241: galois_lookup_251 = 8'hF7;
        8'd242: galois_lookup_251 = 8'h39;
        8'd243: galois_lookup_251 = 8'hC2;
        8'd244: galois_lookup_251 = 8'h66;
        8'd245: galois_lookup_251 = 8'h9D;
        8'd246: galois_lookup_251 = 8'h53;
        8'd247: galois_lookup_251 = 8'hA8;
        8'd248: galois_lookup_251 = 8'hD8;
        8'd249: galois_lookup_251 = 8'h23;
        8'd250: galois_lookup_251 = 8'hED;
        8'd251: galois_lookup_251 = 8'h16;
        8'd252: galois_lookup_251 = 8'hB2;
        8'd253: galois_lookup_251 = 8'h49;
        8'd254: galois_lookup_251 = 8'h87;
        8'd255: galois_lookup_251 = 8'h7C;
    endcase end
endfunction

endmodule

// `endif // LOOKUPS_V
